dff_pre_simulation
.include TSMC_180nm.txt
.include sub_circuits.sub
.include dff.sub

.param LAMBDA=0.09u
.param SUPPLY=1.8
.param width=1.8u

.global vdd gnd

VDD vdd gnd 'SUPPLY'

Vclk clk gnd pulse (1.8 0 0 0 0 5n 10n)

Vd d gnd pulse (0 1.8 3n 0 0 10n 20n) 

Xdff1 q d clk vdd gnd dff

.tran 0.01n 20n

* Measuring tpcq
.measure tran tpcq_r trig v(clk) val='SUPPLY/2' rise=1 targ v(q) val='SUPPLY/2' rise=1
.measure tran tpcq_f trig v(clk) val='SUPPLY/2' rise=2 targ v(q) val='SUPPLY/2' fall=1
.measure tran tpcq param='(tpcq_r+tpcq_f)/2' goal=1

.control
set hcopypscolor = 1 
set color0=white 
set color1=black 

run
set curplottitle=Vedant_Tejas-2023112018-q3-dff
plot v(q) v(d)+2 v(clk)+4
.endc