magic
tech scmos
timestamp 1732087454
<< nwell >>
rect -376 -282 -324 -258
rect -289 -282 -265 -230
rect -376 -322 -324 -298
rect -877 -404 -853 -352
rect -840 -404 -816 -352
rect -921 -451 -895 -411
rect -902 -517 -850 -493
rect -815 -517 -791 -465
rect -532 -486 -508 -434
rect -495 -486 -471 -434
rect -902 -557 -850 -533
rect -680 -548 -656 -496
rect -643 -548 -619 -496
rect -576 -533 -550 -493
rect -366 -536 -314 -512
rect -279 -536 -255 -484
rect -724 -595 -698 -555
rect -366 -576 -314 -552
rect -885 -676 -861 -624
rect -848 -676 -824 -624
rect -929 -723 -903 -683
rect -540 -758 -516 -706
rect -503 -758 -479 -706
rect -910 -841 -858 -817
rect -823 -841 -799 -789
rect -688 -820 -664 -768
rect -651 -820 -627 -768
rect -584 -805 -558 -765
rect -344 -773 -320 -721
rect -307 -773 -283 -721
rect -388 -820 -362 -780
rect -179 -808 -127 -784
rect -92 -808 -68 -756
rect -910 -881 -858 -857
rect -732 -867 -706 -827
rect -179 -848 -127 -824
rect -688 -936 -664 -884
rect -651 -936 -627 -884
rect -732 -983 -706 -943
rect -527 -946 -503 -894
rect -490 -946 -466 -894
rect -571 -993 -545 -953
rect -886 -1107 -862 -1055
rect -849 -1107 -825 -1055
rect -930 -1154 -904 -1114
rect -541 -1189 -517 -1137
rect -504 -1189 -480 -1137
rect -911 -1271 -859 -1247
rect -824 -1271 -800 -1219
rect -689 -1251 -665 -1199
rect -652 -1251 -628 -1199
rect -585 -1236 -559 -1196
rect -345 -1204 -321 -1152
rect -308 -1204 -284 -1152
rect -389 -1251 -363 -1211
rect -180 -1239 -128 -1215
rect -93 -1239 -69 -1187
rect -911 -1311 -859 -1287
rect -733 -1298 -707 -1258
rect -491 -1304 -467 -1252
rect -454 -1304 -430 -1252
rect -180 -1279 -128 -1255
rect -535 -1351 -509 -1311
rect -851 -1410 -827 -1358
rect -814 -1410 -790 -1358
rect -895 -1457 -869 -1417
rect -690 -1420 -666 -1368
rect -653 -1420 -629 -1368
rect -734 -1467 -708 -1427
rect -787 -1605 -763 -1553
rect -750 -1605 -726 -1553
rect -831 -1652 -805 -1612
rect -626 -1615 -602 -1563
rect -589 -1615 -565 -1563
rect -670 -1662 -644 -1622
rect -786 -1723 -762 -1671
rect -749 -1723 -725 -1671
rect -830 -1770 -804 -1730
rect -948 -1859 -924 -1807
rect -911 -1859 -887 -1807
rect -992 -1906 -966 -1866
rect -973 -1972 -921 -1948
rect -886 -1972 -862 -1920
rect -755 -1973 -731 -1921
rect -718 -1973 -694 -1921
rect -603 -1941 -579 -1889
rect -566 -1941 -542 -1889
rect -973 -2012 -921 -1988
rect -799 -2020 -773 -1980
rect -647 -1988 -621 -1948
rect -428 -1972 -404 -1920
rect -391 -1972 -367 -1920
rect -472 -2013 -446 -1979
rect -707 -2158 -683 -2106
rect -670 -2158 -646 -2106
rect -565 -2131 -541 -2079
rect -528 -2131 -504 -2079
rect -751 -2205 -725 -2165
rect -609 -2178 -583 -2138
rect -1076 -2265 -1052 -2213
rect -1039 -2265 -1015 -2213
rect -1120 -2312 -1094 -2272
rect -915 -2275 -891 -2223
rect -878 -2275 -854 -2223
rect -959 -2322 -933 -2282
rect -1021 -2397 -997 -2345
rect -984 -2397 -960 -2345
rect -1065 -2444 -1039 -2404
rect -860 -2407 -836 -2355
rect -823 -2407 -799 -2355
rect -904 -2454 -878 -2414
rect -1020 -2515 -996 -2463
rect -983 -2515 -959 -2463
rect -1064 -2562 -1038 -2522
rect -819 -2644 -795 -2592
rect -782 -2644 -758 -2592
rect -863 -2691 -837 -2651
rect -694 -2675 -670 -2623
rect -657 -2675 -633 -2623
rect -1002 -2771 -978 -2719
rect -965 -2771 -941 -2719
rect -738 -2722 -712 -2682
rect -1046 -2818 -1020 -2778
rect -841 -2781 -817 -2729
rect -804 -2781 -780 -2729
rect -885 -2828 -859 -2788
<< ntransistor >>
rect -404 -271 -384 -269
rect -303 -279 -301 -259
rect -404 -311 -384 -309
rect -303 -317 -301 -297
rect -278 -310 -276 -290
rect -909 -402 -907 -382
rect -866 -432 -864 -412
rect -829 -432 -827 -412
rect -930 -506 -910 -504
rect -829 -514 -827 -494
rect -564 -484 -562 -464
rect -930 -546 -910 -544
rect -829 -552 -827 -532
rect -804 -545 -802 -525
rect -712 -546 -710 -526
rect -521 -514 -519 -494
rect -484 -514 -482 -494
rect -394 -525 -374 -523
rect -293 -533 -291 -513
rect -669 -576 -667 -556
rect -632 -576 -630 -556
rect -394 -565 -374 -563
rect -293 -571 -291 -551
rect -268 -564 -266 -544
rect -917 -674 -915 -654
rect -874 -704 -872 -684
rect -837 -704 -835 -684
rect -572 -756 -570 -736
rect -938 -830 -918 -828
rect -837 -838 -835 -818
rect -720 -818 -718 -798
rect -529 -786 -527 -766
rect -492 -786 -490 -766
rect -376 -771 -374 -751
rect -333 -801 -331 -781
rect -296 -801 -294 -781
rect -207 -797 -187 -795
rect -106 -805 -104 -785
rect -938 -870 -918 -868
rect -837 -876 -835 -856
rect -812 -869 -810 -849
rect -677 -848 -675 -828
rect -640 -848 -638 -828
rect -207 -837 -187 -835
rect -106 -843 -104 -823
rect -81 -836 -79 -816
rect -720 -934 -718 -914
rect -559 -944 -557 -924
rect -677 -964 -675 -944
rect -640 -964 -638 -944
rect -516 -974 -514 -954
rect -479 -974 -477 -954
rect -918 -1105 -916 -1085
rect -875 -1135 -873 -1115
rect -838 -1135 -836 -1115
rect -573 -1187 -571 -1167
rect -939 -1260 -919 -1258
rect -838 -1268 -836 -1248
rect -721 -1249 -719 -1229
rect -530 -1217 -528 -1197
rect -493 -1217 -491 -1197
rect -377 -1202 -375 -1182
rect -334 -1232 -332 -1212
rect -297 -1232 -295 -1212
rect -208 -1228 -188 -1226
rect -107 -1236 -105 -1216
rect -939 -1300 -919 -1298
rect -838 -1306 -836 -1286
rect -813 -1299 -811 -1279
rect -678 -1279 -676 -1259
rect -641 -1279 -639 -1259
rect -523 -1302 -521 -1282
rect -208 -1268 -188 -1266
rect -107 -1274 -105 -1254
rect -82 -1267 -80 -1247
rect -480 -1332 -478 -1312
rect -443 -1332 -441 -1312
rect -883 -1408 -881 -1388
rect -722 -1418 -720 -1398
rect -840 -1438 -838 -1418
rect -803 -1438 -801 -1418
rect -679 -1448 -677 -1428
rect -642 -1448 -640 -1428
rect -819 -1603 -817 -1583
rect -658 -1613 -656 -1593
rect -776 -1633 -774 -1613
rect -739 -1633 -737 -1613
rect -615 -1643 -613 -1623
rect -578 -1643 -576 -1623
rect -818 -1721 -816 -1701
rect -775 -1751 -773 -1731
rect -738 -1751 -736 -1731
rect -980 -1857 -978 -1837
rect -937 -1887 -935 -1867
rect -900 -1887 -898 -1867
rect -1001 -1961 -981 -1959
rect -900 -1969 -898 -1949
rect -787 -1971 -785 -1951
rect -635 -1939 -633 -1919
rect -1001 -2001 -981 -1999
rect -900 -2007 -898 -1987
rect -875 -2000 -873 -1980
rect -592 -1969 -590 -1949
rect -555 -1969 -553 -1949
rect -460 -1970 -458 -1950
rect -744 -2001 -742 -1981
rect -707 -2001 -705 -1981
rect -417 -2000 -415 -1980
rect -380 -2000 -378 -1980
rect -739 -2156 -737 -2136
rect -597 -2129 -595 -2109
rect -554 -2159 -552 -2139
rect -517 -2159 -515 -2139
rect -696 -2186 -694 -2166
rect -659 -2186 -657 -2166
rect -1108 -2263 -1106 -2243
rect -947 -2273 -945 -2253
rect -1065 -2293 -1063 -2273
rect -1028 -2293 -1026 -2273
rect -904 -2303 -902 -2283
rect -867 -2303 -865 -2283
rect -1053 -2395 -1051 -2375
rect -892 -2405 -890 -2385
rect -1010 -2425 -1008 -2405
rect -973 -2425 -971 -2405
rect -849 -2435 -847 -2415
rect -812 -2435 -810 -2415
rect -1052 -2513 -1050 -2493
rect -1009 -2543 -1007 -2523
rect -972 -2543 -970 -2523
rect -851 -2642 -849 -2622
rect -808 -2672 -806 -2652
rect -771 -2672 -769 -2652
rect -726 -2673 -724 -2653
rect -683 -2703 -681 -2683
rect -646 -2703 -644 -2683
rect -1034 -2769 -1032 -2749
rect -873 -2779 -871 -2759
rect -991 -2799 -989 -2779
rect -954 -2799 -952 -2779
rect -830 -2809 -828 -2789
rect -793 -2809 -791 -2789
<< ptransistor >>
rect -370 -271 -330 -269
rect -278 -276 -276 -236
rect -370 -311 -330 -309
rect -866 -398 -864 -358
rect -829 -398 -827 -358
rect -909 -439 -907 -419
rect -896 -506 -856 -504
rect -804 -511 -802 -471
rect -521 -480 -519 -440
rect -484 -480 -482 -440
rect -896 -546 -856 -544
rect -669 -542 -667 -502
rect -632 -542 -630 -502
rect -564 -521 -562 -501
rect -360 -525 -320 -523
rect -268 -530 -266 -490
rect -712 -583 -710 -563
rect -360 -565 -320 -563
rect -874 -670 -872 -630
rect -837 -670 -835 -630
rect -917 -711 -915 -691
rect -529 -752 -527 -712
rect -492 -752 -490 -712
rect -904 -830 -864 -828
rect -812 -835 -810 -795
rect -677 -814 -675 -774
rect -640 -814 -638 -774
rect -572 -793 -570 -773
rect -333 -767 -331 -727
rect -296 -767 -294 -727
rect -376 -808 -374 -788
rect -173 -797 -133 -795
rect -81 -802 -79 -762
rect -904 -870 -864 -868
rect -720 -855 -718 -835
rect -173 -837 -133 -835
rect -677 -930 -675 -890
rect -640 -930 -638 -890
rect -516 -940 -514 -900
rect -479 -940 -477 -900
rect -720 -971 -718 -951
rect -559 -981 -557 -961
rect -875 -1101 -873 -1061
rect -838 -1101 -836 -1061
rect -918 -1142 -916 -1122
rect -530 -1183 -528 -1143
rect -493 -1183 -491 -1143
rect -905 -1260 -865 -1258
rect -813 -1265 -811 -1225
rect -678 -1245 -676 -1205
rect -641 -1245 -639 -1205
rect -573 -1224 -571 -1204
rect -334 -1198 -332 -1158
rect -297 -1198 -295 -1158
rect -377 -1239 -375 -1219
rect -174 -1228 -134 -1226
rect -82 -1233 -80 -1193
rect -905 -1300 -865 -1298
rect -721 -1286 -719 -1266
rect -480 -1298 -478 -1258
rect -443 -1298 -441 -1258
rect -174 -1268 -134 -1266
rect -523 -1339 -521 -1319
rect -840 -1404 -838 -1364
rect -803 -1404 -801 -1364
rect -679 -1414 -677 -1374
rect -642 -1414 -640 -1374
rect -883 -1445 -881 -1425
rect -722 -1455 -720 -1435
rect -776 -1599 -774 -1559
rect -739 -1599 -737 -1559
rect -615 -1609 -613 -1569
rect -578 -1609 -576 -1569
rect -819 -1640 -817 -1620
rect -658 -1650 -656 -1630
rect -775 -1717 -773 -1677
rect -738 -1717 -736 -1677
rect -818 -1758 -816 -1738
rect -937 -1853 -935 -1813
rect -900 -1853 -898 -1813
rect -980 -1894 -978 -1874
rect -967 -1961 -927 -1959
rect -875 -1966 -873 -1926
rect -744 -1967 -742 -1927
rect -707 -1967 -705 -1927
rect -592 -1935 -590 -1895
rect -555 -1935 -553 -1895
rect -967 -2001 -927 -1999
rect -635 -1976 -633 -1956
rect -417 -1966 -415 -1926
rect -380 -1966 -378 -1926
rect -787 -2008 -785 -1988
rect -460 -2007 -458 -1987
rect -696 -2152 -694 -2112
rect -659 -2152 -657 -2112
rect -554 -2125 -552 -2085
rect -517 -2125 -515 -2085
rect -597 -2166 -595 -2146
rect -739 -2193 -737 -2173
rect -1065 -2259 -1063 -2219
rect -1028 -2259 -1026 -2219
rect -904 -2269 -902 -2229
rect -867 -2269 -865 -2229
rect -1108 -2300 -1106 -2280
rect -947 -2310 -945 -2290
rect -1010 -2391 -1008 -2351
rect -973 -2391 -971 -2351
rect -849 -2401 -847 -2361
rect -812 -2401 -810 -2361
rect -1053 -2432 -1051 -2412
rect -892 -2442 -890 -2422
rect -1009 -2509 -1007 -2469
rect -972 -2509 -970 -2469
rect -1052 -2550 -1050 -2530
rect -808 -2638 -806 -2598
rect -771 -2638 -769 -2598
rect -851 -2679 -849 -2659
rect -683 -2669 -681 -2629
rect -646 -2669 -644 -2629
rect -726 -2710 -724 -2690
rect -991 -2765 -989 -2725
rect -954 -2765 -952 -2725
rect -830 -2775 -828 -2735
rect -793 -2775 -791 -2735
rect -1034 -2806 -1032 -2786
rect -873 -2816 -871 -2796
<< ndiffusion >>
rect -404 -269 -384 -268
rect -404 -272 -384 -271
rect -304 -279 -303 -259
rect -301 -279 -300 -259
rect -404 -309 -384 -308
rect -404 -312 -384 -311
rect -304 -317 -303 -297
rect -301 -317 -300 -297
rect -279 -310 -278 -290
rect -276 -310 -275 -290
rect -910 -402 -909 -382
rect -907 -402 -906 -382
rect -867 -432 -866 -412
rect -864 -432 -863 -412
rect -830 -432 -829 -412
rect -827 -432 -826 -412
rect -930 -504 -910 -503
rect -930 -507 -910 -506
rect -830 -514 -829 -494
rect -827 -514 -826 -494
rect -565 -484 -564 -464
rect -562 -484 -561 -464
rect -930 -544 -910 -543
rect -930 -547 -910 -546
rect -830 -552 -829 -532
rect -827 -552 -826 -532
rect -805 -545 -804 -525
rect -802 -545 -801 -525
rect -713 -546 -712 -526
rect -710 -546 -709 -526
rect -522 -514 -521 -494
rect -519 -514 -518 -494
rect -485 -514 -484 -494
rect -482 -514 -481 -494
rect -394 -523 -374 -522
rect -394 -526 -374 -525
rect -294 -533 -293 -513
rect -291 -533 -290 -513
rect -670 -576 -669 -556
rect -667 -576 -666 -556
rect -633 -576 -632 -556
rect -630 -576 -629 -556
rect -394 -563 -374 -562
rect -394 -566 -374 -565
rect -294 -571 -293 -551
rect -291 -571 -290 -551
rect -269 -564 -268 -544
rect -266 -564 -265 -544
rect -918 -674 -917 -654
rect -915 -674 -914 -654
rect -875 -704 -874 -684
rect -872 -704 -871 -684
rect -838 -704 -837 -684
rect -835 -704 -834 -684
rect -573 -756 -572 -736
rect -570 -756 -569 -736
rect -938 -828 -918 -827
rect -938 -831 -918 -830
rect -838 -838 -837 -818
rect -835 -838 -834 -818
rect -721 -818 -720 -798
rect -718 -818 -717 -798
rect -530 -786 -529 -766
rect -527 -786 -526 -766
rect -493 -786 -492 -766
rect -490 -786 -489 -766
rect -377 -771 -376 -751
rect -374 -771 -373 -751
rect -334 -801 -333 -781
rect -331 -801 -330 -781
rect -297 -801 -296 -781
rect -294 -801 -293 -781
rect -207 -795 -187 -794
rect -207 -798 -187 -797
rect -107 -805 -106 -785
rect -104 -805 -103 -785
rect -938 -868 -918 -867
rect -938 -871 -918 -870
rect -838 -876 -837 -856
rect -835 -876 -834 -856
rect -813 -869 -812 -849
rect -810 -869 -809 -849
rect -678 -848 -677 -828
rect -675 -848 -674 -828
rect -641 -848 -640 -828
rect -638 -848 -637 -828
rect -207 -835 -187 -834
rect -207 -838 -187 -837
rect -107 -843 -106 -823
rect -104 -843 -103 -823
rect -82 -836 -81 -816
rect -79 -836 -78 -816
rect -721 -934 -720 -914
rect -718 -934 -717 -914
rect -560 -944 -559 -924
rect -557 -944 -556 -924
rect -678 -964 -677 -944
rect -675 -964 -674 -944
rect -641 -964 -640 -944
rect -638 -964 -637 -944
rect -517 -974 -516 -954
rect -514 -974 -513 -954
rect -480 -974 -479 -954
rect -477 -974 -476 -954
rect -919 -1105 -918 -1085
rect -916 -1105 -915 -1085
rect -876 -1135 -875 -1115
rect -873 -1135 -872 -1115
rect -839 -1135 -838 -1115
rect -836 -1135 -835 -1115
rect -574 -1187 -573 -1167
rect -571 -1187 -570 -1167
rect -939 -1258 -919 -1257
rect -939 -1261 -919 -1260
rect -839 -1268 -838 -1248
rect -836 -1268 -835 -1248
rect -722 -1249 -721 -1229
rect -719 -1249 -718 -1229
rect -531 -1217 -530 -1197
rect -528 -1217 -527 -1197
rect -494 -1217 -493 -1197
rect -491 -1217 -490 -1197
rect -378 -1202 -377 -1182
rect -375 -1202 -374 -1182
rect -335 -1232 -334 -1212
rect -332 -1232 -331 -1212
rect -298 -1232 -297 -1212
rect -295 -1232 -294 -1212
rect -208 -1226 -188 -1225
rect -208 -1229 -188 -1228
rect -108 -1236 -107 -1216
rect -105 -1236 -104 -1216
rect -939 -1298 -919 -1297
rect -939 -1301 -919 -1300
rect -839 -1306 -838 -1286
rect -836 -1306 -835 -1286
rect -814 -1299 -813 -1279
rect -811 -1299 -810 -1279
rect -679 -1279 -678 -1259
rect -676 -1279 -675 -1259
rect -642 -1279 -641 -1259
rect -639 -1279 -638 -1259
rect -524 -1302 -523 -1282
rect -521 -1302 -520 -1282
rect -208 -1266 -188 -1265
rect -208 -1269 -188 -1268
rect -108 -1274 -107 -1254
rect -105 -1274 -104 -1254
rect -83 -1267 -82 -1247
rect -80 -1267 -79 -1247
rect -481 -1332 -480 -1312
rect -478 -1332 -477 -1312
rect -444 -1332 -443 -1312
rect -441 -1332 -440 -1312
rect -884 -1408 -883 -1388
rect -881 -1408 -880 -1388
rect -723 -1418 -722 -1398
rect -720 -1418 -719 -1398
rect -841 -1438 -840 -1418
rect -838 -1438 -837 -1418
rect -804 -1438 -803 -1418
rect -801 -1438 -800 -1418
rect -680 -1448 -679 -1428
rect -677 -1448 -676 -1428
rect -643 -1448 -642 -1428
rect -640 -1448 -639 -1428
rect -820 -1603 -819 -1583
rect -817 -1603 -816 -1583
rect -659 -1613 -658 -1593
rect -656 -1613 -655 -1593
rect -777 -1633 -776 -1613
rect -774 -1633 -773 -1613
rect -740 -1633 -739 -1613
rect -737 -1633 -736 -1613
rect -616 -1643 -615 -1623
rect -613 -1643 -612 -1623
rect -579 -1643 -578 -1623
rect -576 -1643 -575 -1623
rect -819 -1721 -818 -1701
rect -816 -1721 -815 -1701
rect -776 -1751 -775 -1731
rect -773 -1751 -772 -1731
rect -739 -1751 -738 -1731
rect -736 -1751 -735 -1731
rect -981 -1857 -980 -1837
rect -978 -1857 -977 -1837
rect -938 -1887 -937 -1867
rect -935 -1887 -934 -1867
rect -901 -1887 -900 -1867
rect -898 -1887 -897 -1867
rect -1001 -1959 -981 -1958
rect -1001 -1962 -981 -1961
rect -901 -1969 -900 -1949
rect -898 -1969 -897 -1949
rect -788 -1971 -787 -1951
rect -785 -1971 -784 -1951
rect -636 -1939 -635 -1919
rect -633 -1939 -632 -1919
rect -1001 -1999 -981 -1998
rect -1001 -2002 -981 -2001
rect -901 -2007 -900 -1987
rect -898 -2007 -897 -1987
rect -876 -2000 -875 -1980
rect -873 -2000 -872 -1980
rect -593 -1969 -592 -1949
rect -590 -1969 -589 -1949
rect -556 -1969 -555 -1949
rect -553 -1969 -552 -1949
rect -461 -1970 -460 -1950
rect -458 -1970 -457 -1950
rect -745 -2001 -744 -1981
rect -742 -2001 -741 -1981
rect -708 -2001 -707 -1981
rect -705 -2001 -704 -1981
rect -418 -2000 -417 -1980
rect -415 -2000 -414 -1980
rect -381 -2000 -380 -1980
rect -378 -2000 -377 -1980
rect -740 -2156 -739 -2136
rect -737 -2156 -736 -2136
rect -598 -2129 -597 -2109
rect -595 -2129 -594 -2109
rect -555 -2159 -554 -2139
rect -552 -2159 -551 -2139
rect -518 -2159 -517 -2139
rect -515 -2159 -514 -2139
rect -697 -2186 -696 -2166
rect -694 -2186 -693 -2166
rect -660 -2186 -659 -2166
rect -657 -2186 -656 -2166
rect -1109 -2263 -1108 -2243
rect -1106 -2263 -1105 -2243
rect -948 -2273 -947 -2253
rect -945 -2273 -944 -2253
rect -1066 -2293 -1065 -2273
rect -1063 -2293 -1062 -2273
rect -1029 -2293 -1028 -2273
rect -1026 -2293 -1025 -2273
rect -905 -2303 -904 -2283
rect -902 -2303 -901 -2283
rect -868 -2303 -867 -2283
rect -865 -2303 -864 -2283
rect -1054 -2395 -1053 -2375
rect -1051 -2395 -1050 -2375
rect -893 -2405 -892 -2385
rect -890 -2405 -889 -2385
rect -1011 -2425 -1010 -2405
rect -1008 -2425 -1007 -2405
rect -974 -2425 -973 -2405
rect -971 -2425 -970 -2405
rect -850 -2435 -849 -2415
rect -847 -2435 -846 -2415
rect -813 -2435 -812 -2415
rect -810 -2435 -809 -2415
rect -1053 -2513 -1052 -2493
rect -1050 -2513 -1049 -2493
rect -1010 -2543 -1009 -2523
rect -1007 -2543 -1006 -2523
rect -973 -2543 -972 -2523
rect -970 -2543 -969 -2523
rect -852 -2642 -851 -2622
rect -849 -2642 -848 -2622
rect -809 -2672 -808 -2652
rect -806 -2672 -805 -2652
rect -772 -2672 -771 -2652
rect -769 -2672 -768 -2652
rect -727 -2673 -726 -2653
rect -724 -2673 -723 -2653
rect -684 -2703 -683 -2683
rect -681 -2703 -680 -2683
rect -647 -2703 -646 -2683
rect -644 -2703 -643 -2683
rect -1035 -2769 -1034 -2749
rect -1032 -2769 -1031 -2749
rect -874 -2779 -873 -2759
rect -871 -2779 -870 -2759
rect -992 -2799 -991 -2779
rect -989 -2799 -988 -2779
rect -955 -2799 -954 -2779
rect -952 -2799 -951 -2779
rect -831 -2809 -830 -2789
rect -828 -2809 -827 -2789
rect -794 -2809 -793 -2789
rect -791 -2809 -790 -2789
<< pdiffusion >>
rect -370 -269 -330 -268
rect -370 -272 -330 -271
rect -279 -276 -278 -236
rect -276 -276 -275 -236
rect -370 -309 -330 -308
rect -370 -312 -330 -311
rect -867 -398 -866 -358
rect -864 -398 -863 -358
rect -830 -398 -829 -358
rect -827 -398 -826 -358
rect -910 -439 -909 -419
rect -907 -439 -906 -419
rect -896 -504 -856 -503
rect -896 -507 -856 -506
rect -805 -511 -804 -471
rect -802 -511 -801 -471
rect -522 -480 -521 -440
rect -519 -480 -518 -440
rect -485 -480 -484 -440
rect -482 -480 -481 -440
rect -896 -544 -856 -543
rect -896 -547 -856 -546
rect -670 -542 -669 -502
rect -667 -542 -666 -502
rect -633 -542 -632 -502
rect -630 -542 -629 -502
rect -565 -521 -564 -501
rect -562 -521 -561 -501
rect -360 -523 -320 -522
rect -360 -526 -320 -525
rect -269 -530 -268 -490
rect -266 -530 -265 -490
rect -713 -583 -712 -563
rect -710 -583 -709 -563
rect -360 -563 -320 -562
rect -360 -566 -320 -565
rect -875 -670 -874 -630
rect -872 -670 -871 -630
rect -838 -670 -837 -630
rect -835 -670 -834 -630
rect -918 -711 -917 -691
rect -915 -711 -914 -691
rect -530 -752 -529 -712
rect -527 -752 -526 -712
rect -493 -752 -492 -712
rect -490 -752 -489 -712
rect -904 -828 -864 -827
rect -904 -831 -864 -830
rect -813 -835 -812 -795
rect -810 -835 -809 -795
rect -678 -814 -677 -774
rect -675 -814 -674 -774
rect -641 -814 -640 -774
rect -638 -814 -637 -774
rect -573 -793 -572 -773
rect -570 -793 -569 -773
rect -334 -767 -333 -727
rect -331 -767 -330 -727
rect -297 -767 -296 -727
rect -294 -767 -293 -727
rect -377 -808 -376 -788
rect -374 -808 -373 -788
rect -173 -795 -133 -794
rect -173 -798 -133 -797
rect -82 -802 -81 -762
rect -79 -802 -78 -762
rect -904 -868 -864 -867
rect -904 -871 -864 -870
rect -721 -855 -720 -835
rect -718 -855 -717 -835
rect -173 -835 -133 -834
rect -173 -838 -133 -837
rect -678 -930 -677 -890
rect -675 -930 -674 -890
rect -641 -930 -640 -890
rect -638 -930 -637 -890
rect -517 -940 -516 -900
rect -514 -940 -513 -900
rect -480 -940 -479 -900
rect -477 -940 -476 -900
rect -721 -971 -720 -951
rect -718 -971 -717 -951
rect -560 -981 -559 -961
rect -557 -981 -556 -961
rect -876 -1101 -875 -1061
rect -873 -1101 -872 -1061
rect -839 -1101 -838 -1061
rect -836 -1101 -835 -1061
rect -919 -1142 -918 -1122
rect -916 -1142 -915 -1122
rect -531 -1183 -530 -1143
rect -528 -1183 -527 -1143
rect -494 -1183 -493 -1143
rect -491 -1183 -490 -1143
rect -905 -1258 -865 -1257
rect -905 -1261 -865 -1260
rect -814 -1265 -813 -1225
rect -811 -1265 -810 -1225
rect -679 -1245 -678 -1205
rect -676 -1245 -675 -1205
rect -642 -1245 -641 -1205
rect -639 -1245 -638 -1205
rect -574 -1224 -573 -1204
rect -571 -1224 -570 -1204
rect -335 -1198 -334 -1158
rect -332 -1198 -331 -1158
rect -298 -1198 -297 -1158
rect -295 -1198 -294 -1158
rect -378 -1239 -377 -1219
rect -375 -1239 -374 -1219
rect -174 -1226 -134 -1225
rect -174 -1229 -134 -1228
rect -83 -1233 -82 -1193
rect -80 -1233 -79 -1193
rect -905 -1298 -865 -1297
rect -905 -1301 -865 -1300
rect -722 -1286 -721 -1266
rect -719 -1286 -718 -1266
rect -481 -1298 -480 -1258
rect -478 -1298 -477 -1258
rect -444 -1298 -443 -1258
rect -441 -1298 -440 -1258
rect -174 -1266 -134 -1265
rect -174 -1269 -134 -1268
rect -524 -1339 -523 -1319
rect -521 -1339 -520 -1319
rect -841 -1404 -840 -1364
rect -838 -1404 -837 -1364
rect -804 -1404 -803 -1364
rect -801 -1404 -800 -1364
rect -680 -1414 -679 -1374
rect -677 -1414 -676 -1374
rect -643 -1414 -642 -1374
rect -640 -1414 -639 -1374
rect -884 -1445 -883 -1425
rect -881 -1445 -880 -1425
rect -723 -1455 -722 -1435
rect -720 -1455 -719 -1435
rect -777 -1599 -776 -1559
rect -774 -1599 -773 -1559
rect -740 -1599 -739 -1559
rect -737 -1599 -736 -1559
rect -616 -1609 -615 -1569
rect -613 -1609 -612 -1569
rect -579 -1609 -578 -1569
rect -576 -1609 -575 -1569
rect -820 -1640 -819 -1620
rect -817 -1640 -816 -1620
rect -659 -1650 -658 -1630
rect -656 -1650 -655 -1630
rect -776 -1717 -775 -1677
rect -773 -1717 -772 -1677
rect -739 -1717 -738 -1677
rect -736 -1717 -735 -1677
rect -819 -1758 -818 -1738
rect -816 -1758 -815 -1738
rect -938 -1853 -937 -1813
rect -935 -1853 -934 -1813
rect -901 -1853 -900 -1813
rect -898 -1853 -897 -1813
rect -981 -1894 -980 -1874
rect -978 -1894 -977 -1874
rect -967 -1959 -927 -1958
rect -967 -1962 -927 -1961
rect -876 -1966 -875 -1926
rect -873 -1966 -872 -1926
rect -745 -1967 -744 -1927
rect -742 -1967 -741 -1927
rect -708 -1967 -707 -1927
rect -705 -1967 -704 -1927
rect -593 -1935 -592 -1895
rect -590 -1935 -589 -1895
rect -556 -1935 -555 -1895
rect -553 -1935 -552 -1895
rect -967 -1999 -927 -1998
rect -967 -2002 -927 -2001
rect -636 -1976 -635 -1956
rect -633 -1976 -632 -1956
rect -418 -1966 -417 -1926
rect -415 -1966 -414 -1926
rect -381 -1966 -380 -1926
rect -378 -1966 -377 -1926
rect -788 -2008 -787 -1988
rect -785 -2008 -784 -1988
rect -461 -2007 -460 -1987
rect -458 -2007 -457 -1987
rect -697 -2152 -696 -2112
rect -694 -2152 -693 -2112
rect -660 -2152 -659 -2112
rect -657 -2152 -656 -2112
rect -555 -2125 -554 -2085
rect -552 -2125 -551 -2085
rect -518 -2125 -517 -2085
rect -515 -2125 -514 -2085
rect -598 -2166 -597 -2146
rect -595 -2166 -594 -2146
rect -740 -2193 -739 -2173
rect -737 -2193 -736 -2173
rect -1066 -2259 -1065 -2219
rect -1063 -2259 -1062 -2219
rect -1029 -2259 -1028 -2219
rect -1026 -2259 -1025 -2219
rect -905 -2269 -904 -2229
rect -902 -2269 -901 -2229
rect -868 -2269 -867 -2229
rect -865 -2269 -864 -2229
rect -1109 -2300 -1108 -2280
rect -1106 -2300 -1105 -2280
rect -948 -2310 -947 -2290
rect -945 -2310 -944 -2290
rect -1011 -2391 -1010 -2351
rect -1008 -2391 -1007 -2351
rect -974 -2391 -973 -2351
rect -971 -2391 -970 -2351
rect -850 -2401 -849 -2361
rect -847 -2401 -846 -2361
rect -813 -2401 -812 -2361
rect -810 -2401 -809 -2361
rect -1054 -2432 -1053 -2412
rect -1051 -2432 -1050 -2412
rect -893 -2442 -892 -2422
rect -890 -2442 -889 -2422
rect -1010 -2509 -1009 -2469
rect -1007 -2509 -1006 -2469
rect -973 -2509 -972 -2469
rect -970 -2509 -969 -2469
rect -1053 -2550 -1052 -2530
rect -1050 -2550 -1049 -2530
rect -809 -2638 -808 -2598
rect -806 -2638 -805 -2598
rect -772 -2638 -771 -2598
rect -769 -2638 -768 -2598
rect -852 -2679 -851 -2659
rect -849 -2679 -848 -2659
rect -684 -2669 -683 -2629
rect -681 -2669 -680 -2629
rect -647 -2669 -646 -2629
rect -644 -2669 -643 -2629
rect -727 -2710 -726 -2690
rect -724 -2710 -723 -2690
rect -992 -2765 -991 -2725
rect -989 -2765 -988 -2725
rect -955 -2765 -954 -2725
rect -952 -2765 -951 -2725
rect -831 -2775 -830 -2735
rect -828 -2775 -827 -2735
rect -794 -2775 -793 -2735
rect -791 -2775 -790 -2735
rect -1035 -2806 -1034 -2786
rect -1032 -2806 -1031 -2786
rect -874 -2816 -873 -2796
rect -871 -2816 -870 -2796
<< ndcontact >>
rect -404 -268 -384 -264
rect -404 -276 -384 -272
rect -308 -279 -304 -259
rect -300 -279 -296 -259
rect -404 -308 -384 -304
rect -404 -316 -384 -312
rect -308 -317 -304 -297
rect -300 -317 -296 -297
rect -283 -310 -279 -290
rect -275 -310 -271 -290
rect -914 -402 -910 -382
rect -906 -402 -902 -382
rect -871 -432 -867 -412
rect -863 -432 -859 -412
rect -834 -432 -830 -412
rect -826 -432 -822 -412
rect -930 -503 -910 -499
rect -930 -511 -910 -507
rect -834 -514 -830 -494
rect -826 -514 -822 -494
rect -569 -484 -565 -464
rect -561 -484 -557 -464
rect -930 -543 -910 -539
rect -930 -551 -910 -547
rect -834 -552 -830 -532
rect -826 -552 -822 -532
rect -809 -545 -805 -525
rect -801 -545 -797 -525
rect -717 -546 -713 -526
rect -709 -546 -705 -526
rect -526 -514 -522 -494
rect -518 -514 -514 -494
rect -489 -514 -485 -494
rect -481 -514 -477 -494
rect -394 -522 -374 -518
rect -394 -530 -374 -526
rect -298 -533 -294 -513
rect -290 -533 -286 -513
rect -674 -576 -670 -556
rect -666 -576 -662 -556
rect -637 -576 -633 -556
rect -629 -576 -625 -556
rect -394 -562 -374 -558
rect -394 -570 -374 -566
rect -298 -571 -294 -551
rect -290 -571 -286 -551
rect -273 -564 -269 -544
rect -265 -564 -261 -544
rect -922 -674 -918 -654
rect -914 -674 -910 -654
rect -879 -704 -875 -684
rect -871 -704 -867 -684
rect -842 -704 -838 -684
rect -834 -704 -830 -684
rect -577 -756 -573 -736
rect -569 -756 -565 -736
rect -938 -827 -918 -823
rect -938 -835 -918 -831
rect -842 -838 -838 -818
rect -834 -838 -830 -818
rect -725 -818 -721 -798
rect -717 -818 -713 -798
rect -534 -786 -530 -766
rect -526 -786 -522 -766
rect -497 -786 -493 -766
rect -489 -786 -485 -766
rect -381 -771 -377 -751
rect -373 -771 -369 -751
rect -338 -801 -334 -781
rect -330 -801 -326 -781
rect -301 -801 -297 -781
rect -293 -801 -289 -781
rect -207 -794 -187 -790
rect -207 -802 -187 -798
rect -111 -805 -107 -785
rect -103 -805 -99 -785
rect -938 -867 -918 -863
rect -938 -875 -918 -871
rect -842 -876 -838 -856
rect -834 -876 -830 -856
rect -817 -869 -813 -849
rect -809 -869 -805 -849
rect -682 -848 -678 -828
rect -674 -848 -670 -828
rect -645 -848 -641 -828
rect -637 -848 -633 -828
rect -207 -834 -187 -830
rect -207 -842 -187 -838
rect -111 -843 -107 -823
rect -103 -843 -99 -823
rect -86 -836 -82 -816
rect -78 -836 -74 -816
rect -725 -934 -721 -914
rect -717 -934 -713 -914
rect -564 -944 -560 -924
rect -556 -944 -552 -924
rect -682 -964 -678 -944
rect -674 -964 -670 -944
rect -645 -964 -641 -944
rect -637 -964 -633 -944
rect -521 -974 -517 -954
rect -513 -974 -509 -954
rect -484 -974 -480 -954
rect -476 -974 -472 -954
rect -923 -1105 -919 -1085
rect -915 -1105 -911 -1085
rect -880 -1135 -876 -1115
rect -872 -1135 -868 -1115
rect -843 -1135 -839 -1115
rect -835 -1135 -831 -1115
rect -578 -1187 -574 -1167
rect -570 -1187 -566 -1167
rect -939 -1257 -919 -1253
rect -939 -1265 -919 -1261
rect -843 -1268 -839 -1248
rect -835 -1268 -831 -1248
rect -726 -1249 -722 -1229
rect -718 -1249 -714 -1229
rect -535 -1217 -531 -1197
rect -527 -1217 -523 -1197
rect -498 -1217 -494 -1197
rect -490 -1217 -486 -1197
rect -382 -1202 -378 -1182
rect -374 -1202 -370 -1182
rect -339 -1232 -335 -1212
rect -331 -1232 -327 -1212
rect -302 -1232 -298 -1212
rect -294 -1232 -290 -1212
rect -208 -1225 -188 -1221
rect -208 -1233 -188 -1229
rect -112 -1236 -108 -1216
rect -104 -1236 -100 -1216
rect -939 -1297 -919 -1293
rect -939 -1305 -919 -1301
rect -843 -1306 -839 -1286
rect -835 -1306 -831 -1286
rect -818 -1299 -814 -1279
rect -810 -1299 -806 -1279
rect -683 -1279 -679 -1259
rect -675 -1279 -671 -1259
rect -646 -1279 -642 -1259
rect -638 -1279 -634 -1259
rect -528 -1302 -524 -1282
rect -520 -1302 -516 -1282
rect -208 -1265 -188 -1261
rect -208 -1273 -188 -1269
rect -112 -1274 -108 -1254
rect -104 -1274 -100 -1254
rect -87 -1267 -83 -1247
rect -79 -1267 -75 -1247
rect -485 -1332 -481 -1312
rect -477 -1332 -473 -1312
rect -448 -1332 -444 -1312
rect -440 -1332 -436 -1312
rect -888 -1408 -884 -1388
rect -880 -1408 -876 -1388
rect -727 -1418 -723 -1398
rect -719 -1418 -715 -1398
rect -845 -1438 -841 -1418
rect -837 -1438 -833 -1418
rect -808 -1438 -804 -1418
rect -800 -1438 -796 -1418
rect -684 -1448 -680 -1428
rect -676 -1448 -672 -1428
rect -647 -1448 -643 -1428
rect -639 -1448 -635 -1428
rect -824 -1603 -820 -1583
rect -816 -1603 -812 -1583
rect -663 -1613 -659 -1593
rect -655 -1613 -651 -1593
rect -781 -1633 -777 -1613
rect -773 -1633 -769 -1613
rect -744 -1633 -740 -1613
rect -736 -1633 -732 -1613
rect -620 -1643 -616 -1623
rect -612 -1643 -608 -1623
rect -583 -1643 -579 -1623
rect -575 -1643 -571 -1623
rect -823 -1721 -819 -1701
rect -815 -1721 -811 -1701
rect -780 -1751 -776 -1731
rect -772 -1751 -768 -1731
rect -743 -1751 -739 -1731
rect -735 -1751 -731 -1731
rect -985 -1857 -981 -1837
rect -977 -1857 -973 -1837
rect -942 -1887 -938 -1867
rect -934 -1887 -930 -1867
rect -905 -1887 -901 -1867
rect -897 -1887 -893 -1867
rect -1001 -1958 -981 -1954
rect -1001 -1966 -981 -1962
rect -905 -1969 -901 -1949
rect -897 -1969 -893 -1949
rect -792 -1971 -788 -1951
rect -784 -1971 -780 -1951
rect -640 -1939 -636 -1919
rect -632 -1939 -628 -1919
rect -1001 -1998 -981 -1994
rect -1001 -2006 -981 -2002
rect -905 -2007 -901 -1987
rect -897 -2007 -893 -1987
rect -880 -2000 -876 -1980
rect -872 -2000 -868 -1980
rect -597 -1969 -593 -1949
rect -589 -1969 -585 -1949
rect -560 -1969 -556 -1949
rect -552 -1969 -548 -1949
rect -465 -1970 -461 -1950
rect -457 -1970 -453 -1950
rect -749 -2001 -745 -1981
rect -741 -2001 -737 -1981
rect -712 -2001 -708 -1981
rect -704 -2001 -700 -1981
rect -422 -2000 -418 -1980
rect -414 -2000 -410 -1980
rect -385 -2000 -381 -1980
rect -377 -2000 -373 -1980
rect -744 -2156 -740 -2136
rect -736 -2156 -732 -2136
rect -602 -2129 -598 -2109
rect -594 -2129 -590 -2109
rect -559 -2159 -555 -2139
rect -551 -2159 -547 -2139
rect -522 -2159 -518 -2139
rect -514 -2159 -510 -2139
rect -701 -2186 -697 -2166
rect -693 -2186 -689 -2166
rect -664 -2186 -660 -2166
rect -656 -2186 -652 -2166
rect -1113 -2263 -1109 -2243
rect -1105 -2263 -1101 -2243
rect -952 -2273 -948 -2253
rect -944 -2273 -940 -2253
rect -1070 -2293 -1066 -2273
rect -1062 -2293 -1058 -2273
rect -1033 -2293 -1029 -2273
rect -1025 -2293 -1021 -2273
rect -909 -2303 -905 -2283
rect -901 -2303 -897 -2283
rect -872 -2303 -868 -2283
rect -864 -2303 -860 -2283
rect -1058 -2395 -1054 -2375
rect -1050 -2395 -1046 -2375
rect -897 -2405 -893 -2385
rect -889 -2405 -885 -2385
rect -1015 -2425 -1011 -2405
rect -1007 -2425 -1003 -2405
rect -978 -2425 -974 -2405
rect -970 -2425 -966 -2405
rect -854 -2435 -850 -2415
rect -846 -2435 -842 -2415
rect -817 -2435 -813 -2415
rect -809 -2435 -805 -2415
rect -1057 -2513 -1053 -2493
rect -1049 -2513 -1045 -2493
rect -1014 -2543 -1010 -2523
rect -1006 -2543 -1002 -2523
rect -977 -2543 -973 -2523
rect -969 -2543 -965 -2523
rect -856 -2642 -852 -2622
rect -848 -2642 -844 -2622
rect -813 -2672 -809 -2652
rect -805 -2672 -801 -2652
rect -776 -2672 -772 -2652
rect -768 -2672 -764 -2652
rect -731 -2673 -727 -2653
rect -723 -2673 -719 -2653
rect -688 -2703 -684 -2683
rect -680 -2703 -676 -2683
rect -651 -2703 -647 -2683
rect -643 -2703 -639 -2683
rect -1039 -2769 -1035 -2749
rect -1031 -2769 -1027 -2749
rect -878 -2779 -874 -2759
rect -870 -2779 -866 -2759
rect -996 -2799 -992 -2779
rect -988 -2799 -984 -2779
rect -959 -2799 -955 -2779
rect -951 -2799 -947 -2779
rect -835 -2809 -831 -2789
rect -827 -2809 -823 -2789
rect -798 -2809 -794 -2789
rect -790 -2809 -786 -2789
<< pdcontact >>
rect -370 -268 -330 -264
rect -370 -276 -330 -272
rect -283 -276 -279 -236
rect -275 -276 -271 -236
rect -370 -308 -330 -304
rect -370 -316 -330 -312
rect -871 -398 -867 -358
rect -863 -398 -859 -358
rect -834 -398 -830 -358
rect -826 -398 -822 -358
rect -914 -439 -910 -419
rect -906 -439 -902 -419
rect -896 -503 -856 -499
rect -896 -511 -856 -507
rect -809 -511 -805 -471
rect -801 -511 -797 -471
rect -526 -480 -522 -440
rect -518 -480 -514 -440
rect -489 -480 -485 -440
rect -481 -480 -477 -440
rect -896 -543 -856 -539
rect -896 -551 -856 -547
rect -674 -542 -670 -502
rect -666 -542 -662 -502
rect -637 -542 -633 -502
rect -629 -542 -625 -502
rect -569 -521 -565 -501
rect -561 -521 -557 -501
rect -360 -522 -320 -518
rect -360 -530 -320 -526
rect -273 -530 -269 -490
rect -265 -530 -261 -490
rect -717 -583 -713 -563
rect -709 -583 -705 -563
rect -360 -562 -320 -558
rect -360 -570 -320 -566
rect -879 -670 -875 -630
rect -871 -670 -867 -630
rect -842 -670 -838 -630
rect -834 -670 -830 -630
rect -922 -711 -918 -691
rect -914 -711 -910 -691
rect -534 -752 -530 -712
rect -526 -752 -522 -712
rect -497 -752 -493 -712
rect -489 -752 -485 -712
rect -904 -827 -864 -823
rect -904 -835 -864 -831
rect -817 -835 -813 -795
rect -809 -835 -805 -795
rect -682 -814 -678 -774
rect -674 -814 -670 -774
rect -645 -814 -641 -774
rect -637 -814 -633 -774
rect -577 -793 -573 -773
rect -569 -793 -565 -773
rect -338 -767 -334 -727
rect -330 -767 -326 -727
rect -301 -767 -297 -727
rect -293 -767 -289 -727
rect -381 -808 -377 -788
rect -373 -808 -369 -788
rect -173 -794 -133 -790
rect -173 -802 -133 -798
rect -86 -802 -82 -762
rect -78 -802 -74 -762
rect -904 -867 -864 -863
rect -904 -875 -864 -871
rect -725 -855 -721 -835
rect -717 -855 -713 -835
rect -173 -834 -133 -830
rect -173 -842 -133 -838
rect -682 -930 -678 -890
rect -674 -930 -670 -890
rect -645 -930 -641 -890
rect -637 -930 -633 -890
rect -521 -940 -517 -900
rect -513 -940 -509 -900
rect -484 -940 -480 -900
rect -476 -940 -472 -900
rect -725 -971 -721 -951
rect -717 -971 -713 -951
rect -564 -981 -560 -961
rect -556 -981 -552 -961
rect -880 -1101 -876 -1061
rect -872 -1101 -868 -1061
rect -843 -1101 -839 -1061
rect -835 -1101 -831 -1061
rect -923 -1142 -919 -1122
rect -915 -1142 -911 -1122
rect -535 -1183 -531 -1143
rect -527 -1183 -523 -1143
rect -498 -1183 -494 -1143
rect -490 -1183 -486 -1143
rect -905 -1257 -865 -1253
rect -905 -1265 -865 -1261
rect -818 -1265 -814 -1225
rect -810 -1265 -806 -1225
rect -683 -1245 -679 -1205
rect -675 -1245 -671 -1205
rect -646 -1245 -642 -1205
rect -638 -1245 -634 -1205
rect -578 -1224 -574 -1204
rect -570 -1224 -566 -1204
rect -339 -1198 -335 -1158
rect -331 -1198 -327 -1158
rect -302 -1198 -298 -1158
rect -294 -1198 -290 -1158
rect -382 -1239 -378 -1219
rect -374 -1239 -370 -1219
rect -174 -1225 -134 -1221
rect -174 -1233 -134 -1229
rect -87 -1233 -83 -1193
rect -79 -1233 -75 -1193
rect -905 -1297 -865 -1293
rect -905 -1305 -865 -1301
rect -726 -1286 -722 -1266
rect -718 -1286 -714 -1266
rect -485 -1298 -481 -1258
rect -477 -1298 -473 -1258
rect -448 -1298 -444 -1258
rect -440 -1298 -436 -1258
rect -174 -1265 -134 -1261
rect -174 -1273 -134 -1269
rect -528 -1339 -524 -1319
rect -520 -1339 -516 -1319
rect -845 -1404 -841 -1364
rect -837 -1404 -833 -1364
rect -808 -1404 -804 -1364
rect -800 -1404 -796 -1364
rect -684 -1414 -680 -1374
rect -676 -1414 -672 -1374
rect -647 -1414 -643 -1374
rect -639 -1414 -635 -1374
rect -888 -1445 -884 -1425
rect -880 -1445 -876 -1425
rect -727 -1455 -723 -1435
rect -719 -1455 -715 -1435
rect -781 -1599 -777 -1559
rect -773 -1599 -769 -1559
rect -744 -1599 -740 -1559
rect -736 -1599 -732 -1559
rect -620 -1609 -616 -1569
rect -612 -1609 -608 -1569
rect -583 -1609 -579 -1569
rect -575 -1609 -571 -1569
rect -824 -1640 -820 -1620
rect -816 -1640 -812 -1620
rect -663 -1650 -659 -1630
rect -655 -1650 -651 -1630
rect -780 -1717 -776 -1677
rect -772 -1717 -768 -1677
rect -743 -1717 -739 -1677
rect -735 -1717 -731 -1677
rect -823 -1758 -819 -1738
rect -815 -1758 -811 -1738
rect -942 -1853 -938 -1813
rect -934 -1853 -930 -1813
rect -905 -1853 -901 -1813
rect -897 -1853 -893 -1813
rect -985 -1894 -981 -1874
rect -977 -1894 -973 -1874
rect -967 -1958 -927 -1954
rect -967 -1966 -927 -1962
rect -880 -1966 -876 -1926
rect -872 -1966 -868 -1926
rect -749 -1967 -745 -1927
rect -741 -1967 -737 -1927
rect -712 -1967 -708 -1927
rect -704 -1967 -700 -1927
rect -597 -1935 -593 -1895
rect -589 -1935 -585 -1895
rect -560 -1935 -556 -1895
rect -552 -1935 -548 -1895
rect -967 -1998 -927 -1994
rect -967 -2006 -927 -2002
rect -640 -1976 -636 -1956
rect -632 -1976 -628 -1956
rect -422 -1966 -418 -1926
rect -414 -1966 -410 -1926
rect -385 -1966 -381 -1926
rect -377 -1966 -373 -1926
rect -792 -2008 -788 -1988
rect -784 -2008 -780 -1988
rect -465 -2007 -461 -1987
rect -457 -2007 -453 -1987
rect -701 -2152 -697 -2112
rect -693 -2152 -689 -2112
rect -664 -2152 -660 -2112
rect -656 -2152 -652 -2112
rect -559 -2125 -555 -2085
rect -551 -2125 -547 -2085
rect -522 -2125 -518 -2085
rect -514 -2125 -510 -2085
rect -602 -2166 -598 -2146
rect -594 -2166 -590 -2146
rect -744 -2193 -740 -2173
rect -736 -2193 -732 -2173
rect -1070 -2259 -1066 -2219
rect -1062 -2259 -1058 -2219
rect -1033 -2259 -1029 -2219
rect -1025 -2259 -1021 -2219
rect -909 -2269 -905 -2229
rect -901 -2269 -897 -2229
rect -872 -2269 -868 -2229
rect -864 -2269 -860 -2229
rect -1113 -2300 -1109 -2280
rect -1105 -2300 -1101 -2280
rect -952 -2310 -948 -2290
rect -944 -2310 -940 -2290
rect -1015 -2391 -1011 -2351
rect -1007 -2391 -1003 -2351
rect -978 -2391 -974 -2351
rect -970 -2391 -966 -2351
rect -854 -2401 -850 -2361
rect -846 -2401 -842 -2361
rect -817 -2401 -813 -2361
rect -809 -2401 -805 -2361
rect -1058 -2432 -1054 -2412
rect -1050 -2432 -1046 -2412
rect -897 -2442 -893 -2422
rect -889 -2442 -885 -2422
rect -1014 -2509 -1010 -2469
rect -1006 -2509 -1002 -2469
rect -977 -2509 -973 -2469
rect -969 -2509 -965 -2469
rect -1057 -2550 -1053 -2530
rect -1049 -2550 -1045 -2530
rect -813 -2638 -809 -2598
rect -805 -2638 -801 -2598
rect -776 -2638 -772 -2598
rect -768 -2638 -764 -2598
rect -856 -2679 -852 -2659
rect -848 -2679 -844 -2659
rect -688 -2669 -684 -2629
rect -680 -2669 -676 -2629
rect -651 -2669 -647 -2629
rect -643 -2669 -639 -2629
rect -731 -2710 -727 -2690
rect -723 -2710 -719 -2690
rect -996 -2765 -992 -2725
rect -988 -2765 -984 -2725
rect -959 -2765 -955 -2725
rect -951 -2765 -947 -2725
rect -835 -2775 -831 -2735
rect -827 -2775 -823 -2735
rect -798 -2775 -794 -2735
rect -790 -2775 -786 -2735
rect -1039 -2806 -1035 -2786
rect -1031 -2806 -1027 -2786
rect -878 -2816 -874 -2796
rect -870 -2816 -866 -2796
<< psubstratepcontact >>
rect -414 -263 -410 -259
rect -414 -281 -410 -277
rect -414 -303 -410 -299
rect -414 -321 -410 -317
rect -288 -320 -284 -316
rect -270 -320 -266 -316
rect -876 -442 -872 -438
rect -858 -442 -854 -438
rect -839 -442 -835 -438
rect -821 -442 -817 -438
rect -940 -498 -936 -494
rect -940 -516 -936 -512
rect -940 -538 -936 -534
rect -940 -556 -936 -552
rect -404 -517 -400 -513
rect -531 -524 -527 -520
rect -513 -524 -509 -520
rect -494 -524 -490 -520
rect -476 -524 -472 -520
rect -404 -535 -400 -531
rect -814 -555 -810 -551
rect -796 -555 -792 -551
rect -404 -557 -400 -553
rect -404 -575 -400 -571
rect -278 -574 -274 -570
rect -260 -574 -256 -570
rect -679 -586 -675 -582
rect -661 -586 -657 -582
rect -642 -586 -638 -582
rect -624 -586 -620 -582
rect -884 -714 -880 -710
rect -866 -714 -862 -710
rect -847 -714 -843 -710
rect -829 -714 -825 -710
rect -948 -822 -944 -818
rect -948 -840 -944 -836
rect -539 -796 -535 -792
rect -521 -796 -517 -792
rect -502 -796 -498 -792
rect -484 -796 -480 -792
rect -217 -789 -213 -785
rect -217 -807 -213 -803
rect -343 -811 -339 -807
rect -325 -811 -321 -807
rect -306 -811 -302 -807
rect -288 -811 -284 -807
rect -948 -862 -944 -858
rect -948 -880 -944 -876
rect -217 -829 -213 -825
rect -217 -847 -213 -843
rect -91 -846 -87 -842
rect -73 -846 -69 -842
rect -687 -858 -683 -854
rect -669 -858 -665 -854
rect -650 -858 -646 -854
rect -632 -858 -628 -854
rect -822 -879 -818 -875
rect -804 -879 -800 -875
rect -687 -974 -683 -970
rect -669 -974 -665 -970
rect -650 -974 -646 -970
rect -632 -974 -628 -970
rect -526 -984 -522 -980
rect -508 -984 -504 -980
rect -489 -984 -485 -980
rect -471 -984 -467 -980
rect -885 -1145 -881 -1141
rect -867 -1145 -863 -1141
rect -848 -1145 -844 -1141
rect -830 -1145 -826 -1141
rect -949 -1252 -945 -1248
rect -949 -1270 -945 -1266
rect -540 -1227 -536 -1223
rect -522 -1227 -518 -1223
rect -503 -1227 -499 -1223
rect -485 -1227 -481 -1223
rect -218 -1220 -214 -1216
rect -218 -1238 -214 -1234
rect -344 -1242 -340 -1238
rect -326 -1242 -322 -1238
rect -307 -1242 -303 -1238
rect -289 -1242 -285 -1238
rect -949 -1292 -945 -1288
rect -949 -1310 -945 -1306
rect -688 -1289 -684 -1285
rect -670 -1289 -666 -1285
rect -651 -1289 -647 -1285
rect -633 -1289 -629 -1285
rect -218 -1260 -214 -1256
rect -218 -1278 -214 -1274
rect -92 -1277 -88 -1273
rect -74 -1277 -70 -1273
rect -823 -1309 -819 -1305
rect -805 -1309 -801 -1305
rect -490 -1342 -486 -1338
rect -472 -1342 -468 -1338
rect -453 -1342 -449 -1338
rect -435 -1342 -431 -1338
rect -850 -1448 -846 -1444
rect -832 -1448 -828 -1444
rect -813 -1448 -809 -1444
rect -795 -1448 -791 -1444
rect -689 -1458 -685 -1454
rect -671 -1458 -667 -1454
rect -652 -1458 -648 -1454
rect -634 -1458 -630 -1454
rect -786 -1643 -782 -1639
rect -768 -1643 -764 -1639
rect -749 -1643 -745 -1639
rect -731 -1643 -727 -1639
rect -625 -1653 -621 -1649
rect -607 -1653 -603 -1649
rect -588 -1653 -584 -1649
rect -570 -1653 -566 -1649
rect -785 -1761 -781 -1757
rect -767 -1761 -763 -1757
rect -748 -1761 -744 -1757
rect -730 -1761 -726 -1757
rect -947 -1897 -943 -1893
rect -929 -1897 -925 -1893
rect -910 -1897 -906 -1893
rect -892 -1897 -888 -1893
rect -1011 -1953 -1007 -1949
rect -1011 -1971 -1007 -1967
rect -1011 -1993 -1007 -1989
rect -1011 -2011 -1007 -2007
rect -602 -1979 -598 -1975
rect -584 -1979 -580 -1975
rect -565 -1979 -561 -1975
rect -547 -1979 -543 -1975
rect -885 -2010 -881 -2006
rect -867 -2010 -863 -2006
rect -754 -2011 -750 -2007
rect -736 -2011 -732 -2007
rect -717 -2011 -713 -2007
rect -699 -2011 -695 -2007
rect -427 -2010 -423 -2006
rect -409 -2010 -405 -2006
rect -390 -2010 -386 -2006
rect -372 -2010 -368 -2006
rect -564 -2169 -560 -2165
rect -546 -2169 -542 -2165
rect -527 -2169 -523 -2165
rect -509 -2169 -505 -2165
rect -706 -2196 -702 -2192
rect -688 -2196 -684 -2192
rect -669 -2196 -665 -2192
rect -651 -2196 -647 -2192
rect -1075 -2303 -1071 -2299
rect -1057 -2303 -1053 -2299
rect -1038 -2303 -1034 -2299
rect -1020 -2303 -1016 -2299
rect -914 -2313 -910 -2309
rect -896 -2313 -892 -2309
rect -877 -2313 -873 -2309
rect -859 -2313 -855 -2309
rect -1020 -2435 -1016 -2431
rect -1002 -2435 -998 -2431
rect -983 -2435 -979 -2431
rect -965 -2435 -961 -2431
rect -859 -2445 -855 -2441
rect -841 -2445 -837 -2441
rect -822 -2445 -818 -2441
rect -804 -2445 -800 -2441
rect -1019 -2553 -1015 -2549
rect -1001 -2553 -997 -2549
rect -982 -2553 -978 -2549
rect -964 -2553 -960 -2549
rect -818 -2682 -814 -2678
rect -800 -2682 -796 -2678
rect -781 -2682 -777 -2678
rect -763 -2682 -759 -2678
rect -693 -2713 -689 -2709
rect -675 -2713 -671 -2709
rect -656 -2713 -652 -2709
rect -638 -2713 -634 -2709
rect -1001 -2809 -997 -2805
rect -983 -2809 -979 -2805
rect -964 -2809 -960 -2805
rect -946 -2809 -942 -2805
rect -840 -2819 -836 -2815
rect -822 -2819 -818 -2815
rect -803 -2819 -799 -2815
rect -785 -2819 -781 -2815
<< nsubstratencontact >>
rect -286 -228 -282 -224
rect -272 -228 -268 -224
rect -322 -265 -318 -261
rect -322 -279 -318 -275
rect -322 -305 -318 -301
rect -322 -319 -318 -315
rect -874 -350 -870 -346
rect -860 -350 -856 -346
rect -837 -350 -833 -346
rect -823 -350 -819 -346
rect -529 -432 -525 -428
rect -515 -432 -511 -428
rect -492 -432 -488 -428
rect -478 -432 -474 -428
rect -812 -463 -808 -459
rect -798 -463 -794 -459
rect -848 -500 -844 -496
rect -848 -514 -844 -510
rect -677 -494 -673 -490
rect -663 -494 -659 -490
rect -640 -494 -636 -490
rect -626 -494 -622 -490
rect -276 -482 -272 -478
rect -262 -482 -258 -478
rect -848 -540 -844 -536
rect -848 -554 -844 -550
rect -312 -519 -308 -515
rect -312 -533 -308 -529
rect -312 -559 -308 -555
rect -312 -573 -308 -569
rect -882 -622 -878 -618
rect -868 -622 -864 -618
rect -845 -622 -841 -618
rect -831 -622 -827 -618
rect -537 -704 -533 -700
rect -523 -704 -519 -700
rect -500 -704 -496 -700
rect -486 -704 -482 -700
rect -341 -719 -337 -715
rect -327 -719 -323 -715
rect -304 -719 -300 -715
rect -290 -719 -286 -715
rect -685 -766 -681 -762
rect -671 -766 -667 -762
rect -648 -766 -644 -762
rect -634 -766 -630 -762
rect -820 -787 -816 -783
rect -806 -787 -802 -783
rect -856 -824 -852 -820
rect -856 -838 -852 -834
rect -89 -754 -85 -750
rect -75 -754 -71 -750
rect -125 -791 -121 -787
rect -125 -805 -121 -801
rect -856 -864 -852 -860
rect -856 -878 -852 -874
rect -125 -831 -121 -827
rect -125 -845 -121 -841
rect -685 -882 -681 -878
rect -671 -882 -667 -878
rect -648 -882 -644 -878
rect -634 -882 -630 -878
rect -524 -892 -520 -888
rect -510 -892 -506 -888
rect -487 -892 -483 -888
rect -473 -892 -469 -888
rect -883 -1053 -879 -1049
rect -869 -1053 -865 -1049
rect -846 -1053 -842 -1049
rect -832 -1053 -828 -1049
rect -538 -1135 -534 -1131
rect -524 -1135 -520 -1131
rect -501 -1135 -497 -1131
rect -487 -1135 -483 -1131
rect -342 -1150 -338 -1146
rect -328 -1150 -324 -1146
rect -305 -1150 -301 -1146
rect -291 -1150 -287 -1146
rect -686 -1197 -682 -1193
rect -672 -1197 -668 -1193
rect -649 -1197 -645 -1193
rect -635 -1197 -631 -1193
rect -821 -1217 -817 -1213
rect -807 -1217 -803 -1213
rect -857 -1254 -853 -1250
rect -857 -1268 -853 -1264
rect -90 -1185 -86 -1181
rect -76 -1185 -72 -1181
rect -126 -1222 -122 -1218
rect -126 -1236 -122 -1232
rect -488 -1250 -484 -1246
rect -474 -1250 -470 -1246
rect -451 -1250 -447 -1246
rect -437 -1250 -433 -1246
rect -857 -1294 -853 -1290
rect -857 -1308 -853 -1304
rect -126 -1262 -122 -1258
rect -126 -1276 -122 -1272
rect -848 -1356 -844 -1352
rect -834 -1356 -830 -1352
rect -811 -1356 -807 -1352
rect -797 -1356 -793 -1352
rect -687 -1366 -683 -1362
rect -673 -1366 -669 -1362
rect -650 -1366 -646 -1362
rect -636 -1366 -632 -1362
rect -784 -1551 -780 -1547
rect -770 -1551 -766 -1547
rect -747 -1551 -743 -1547
rect -733 -1551 -729 -1547
rect -623 -1561 -619 -1557
rect -609 -1561 -605 -1557
rect -586 -1561 -582 -1557
rect -572 -1561 -568 -1557
rect -783 -1669 -779 -1665
rect -769 -1669 -765 -1665
rect -746 -1669 -742 -1665
rect -732 -1669 -728 -1665
rect -945 -1805 -941 -1801
rect -931 -1805 -927 -1801
rect -908 -1805 -904 -1801
rect -894 -1805 -890 -1801
rect -600 -1887 -596 -1883
rect -586 -1887 -582 -1883
rect -563 -1887 -559 -1883
rect -549 -1887 -545 -1883
rect -883 -1918 -879 -1914
rect -869 -1918 -865 -1914
rect -752 -1919 -748 -1915
rect -738 -1919 -734 -1915
rect -715 -1919 -711 -1915
rect -701 -1919 -697 -1915
rect -919 -1955 -915 -1951
rect -919 -1969 -915 -1965
rect -425 -1918 -421 -1914
rect -411 -1918 -407 -1914
rect -388 -1918 -384 -1914
rect -374 -1918 -370 -1914
rect -919 -1995 -915 -1991
rect -919 -2009 -915 -2005
rect -562 -2077 -558 -2073
rect -548 -2077 -544 -2073
rect -525 -2077 -521 -2073
rect -511 -2077 -507 -2073
rect -704 -2104 -700 -2100
rect -690 -2104 -686 -2100
rect -667 -2104 -663 -2100
rect -653 -2104 -649 -2100
rect -1073 -2211 -1069 -2207
rect -1059 -2211 -1055 -2207
rect -1036 -2211 -1032 -2207
rect -1022 -2211 -1018 -2207
rect -912 -2221 -908 -2217
rect -898 -2221 -894 -2217
rect -875 -2221 -871 -2217
rect -861 -2221 -857 -2217
rect -1018 -2343 -1014 -2339
rect -1004 -2343 -1000 -2339
rect -981 -2343 -977 -2339
rect -967 -2343 -963 -2339
rect -857 -2353 -853 -2349
rect -843 -2353 -839 -2349
rect -820 -2353 -816 -2349
rect -806 -2353 -802 -2349
rect -1017 -2461 -1013 -2457
rect -1003 -2461 -999 -2457
rect -980 -2461 -976 -2457
rect -966 -2461 -962 -2457
rect -816 -2590 -812 -2586
rect -802 -2590 -798 -2586
rect -779 -2590 -775 -2586
rect -765 -2590 -761 -2586
rect -691 -2621 -687 -2617
rect -677 -2621 -673 -2617
rect -654 -2621 -650 -2617
rect -640 -2621 -636 -2617
rect -999 -2717 -995 -2713
rect -985 -2717 -981 -2713
rect -962 -2717 -958 -2713
rect -948 -2717 -944 -2713
rect -838 -2727 -834 -2723
rect -824 -2727 -820 -2723
rect -801 -2727 -797 -2723
rect -787 -2727 -783 -2723
<< polysilicon >>
rect -278 -236 -276 -233
rect -381 -248 -301 -246
rect -303 -259 -301 -248
rect -408 -271 -404 -269
rect -384 -271 -370 -269
rect -330 -271 -327 -269
rect -303 -283 -301 -279
rect -381 -288 -301 -286
rect -303 -297 -301 -288
rect -278 -290 -276 -276
rect -408 -311 -404 -309
rect -384 -311 -370 -309
rect -330 -311 -327 -309
rect -278 -314 -276 -310
rect -303 -321 -301 -317
rect -866 -358 -864 -355
rect -829 -358 -827 -355
rect -909 -382 -907 -374
rect -909 -419 -907 -402
rect -866 -412 -864 -398
rect -829 -412 -827 -398
rect -866 -436 -864 -432
rect -829 -436 -827 -432
rect -909 -443 -907 -439
rect -521 -440 -519 -437
rect -484 -440 -482 -437
rect -564 -464 -562 -456
rect -804 -471 -802 -468
rect -907 -483 -827 -481
rect -829 -494 -827 -483
rect -934 -506 -930 -504
rect -910 -506 -896 -504
rect -856 -506 -853 -504
rect -669 -502 -667 -499
rect -632 -502 -630 -499
rect -564 -501 -562 -484
rect -521 -494 -519 -480
rect -484 -494 -482 -480
rect -268 -490 -266 -487
rect -829 -518 -827 -514
rect -907 -523 -827 -521
rect -829 -532 -827 -523
rect -804 -525 -802 -511
rect -934 -546 -930 -544
rect -910 -546 -896 -544
rect -856 -546 -853 -544
rect -712 -526 -710 -518
rect -804 -549 -802 -545
rect -371 -502 -291 -500
rect -293 -513 -291 -502
rect -521 -518 -519 -514
rect -484 -518 -482 -514
rect -564 -525 -562 -521
rect -398 -525 -394 -523
rect -374 -525 -360 -523
rect -320 -525 -317 -523
rect -293 -537 -291 -533
rect -371 -542 -291 -540
rect -829 -556 -827 -552
rect -712 -563 -710 -546
rect -669 -556 -667 -542
rect -632 -556 -630 -542
rect -293 -551 -291 -542
rect -268 -544 -266 -530
rect -398 -565 -394 -563
rect -374 -565 -360 -563
rect -320 -565 -317 -563
rect -268 -568 -266 -564
rect -293 -575 -291 -571
rect -669 -580 -667 -576
rect -632 -580 -630 -576
rect -712 -587 -710 -583
rect -874 -630 -872 -627
rect -837 -630 -835 -627
rect -917 -654 -915 -646
rect -917 -691 -915 -674
rect -874 -684 -872 -670
rect -837 -684 -835 -670
rect -874 -708 -872 -704
rect -837 -708 -835 -704
rect -917 -715 -915 -711
rect -529 -712 -527 -709
rect -492 -712 -490 -709
rect -572 -736 -570 -728
rect -333 -727 -331 -724
rect -296 -727 -294 -724
rect -376 -751 -374 -743
rect -677 -774 -675 -771
rect -640 -774 -638 -771
rect -572 -773 -570 -756
rect -529 -766 -527 -752
rect -492 -766 -490 -752
rect -812 -795 -810 -792
rect -915 -807 -835 -805
rect -837 -818 -835 -807
rect -942 -830 -938 -828
rect -918 -830 -904 -828
rect -864 -830 -861 -828
rect -720 -798 -718 -790
rect -81 -762 -79 -759
rect -529 -790 -527 -786
rect -492 -790 -490 -786
rect -376 -788 -374 -771
rect -333 -781 -331 -767
rect -296 -781 -294 -767
rect -184 -774 -104 -772
rect -572 -797 -570 -793
rect -106 -785 -104 -774
rect -211 -797 -207 -795
rect -187 -797 -173 -795
rect -133 -797 -130 -795
rect -333 -805 -331 -801
rect -296 -805 -294 -801
rect -376 -812 -374 -808
rect -106 -809 -104 -805
rect -184 -814 -104 -812
rect -720 -835 -718 -818
rect -677 -828 -675 -814
rect -640 -828 -638 -814
rect -106 -823 -104 -814
rect -81 -816 -79 -802
rect -837 -842 -835 -838
rect -915 -847 -835 -845
rect -837 -856 -835 -847
rect -812 -849 -810 -835
rect -942 -870 -938 -868
rect -918 -870 -904 -868
rect -864 -870 -861 -868
rect -211 -837 -207 -835
rect -187 -837 -173 -835
rect -133 -837 -130 -835
rect -81 -840 -79 -836
rect -106 -847 -104 -843
rect -677 -852 -675 -848
rect -640 -852 -638 -848
rect -720 -859 -718 -855
rect -812 -873 -810 -869
rect -837 -880 -835 -876
rect -677 -890 -675 -887
rect -640 -890 -638 -887
rect -720 -914 -718 -906
rect -516 -900 -514 -897
rect -479 -900 -477 -897
rect -559 -924 -557 -916
rect -720 -951 -718 -934
rect -677 -944 -675 -930
rect -640 -944 -638 -930
rect -559 -961 -557 -944
rect -516 -954 -514 -940
rect -479 -954 -477 -940
rect -677 -968 -675 -964
rect -640 -968 -638 -964
rect -720 -975 -718 -971
rect -516 -978 -514 -974
rect -479 -978 -477 -974
rect -559 -985 -557 -981
rect -875 -1061 -873 -1058
rect -838 -1061 -836 -1058
rect -918 -1085 -916 -1077
rect -918 -1122 -916 -1105
rect -875 -1115 -873 -1101
rect -838 -1115 -836 -1101
rect -875 -1139 -873 -1135
rect -838 -1139 -836 -1135
rect -918 -1146 -916 -1142
rect -530 -1143 -528 -1140
rect -493 -1143 -491 -1140
rect -573 -1167 -571 -1159
rect -334 -1158 -332 -1155
rect -297 -1158 -295 -1155
rect -377 -1182 -375 -1174
rect -678 -1205 -676 -1202
rect -641 -1205 -639 -1202
rect -573 -1204 -571 -1187
rect -530 -1197 -528 -1183
rect -493 -1197 -491 -1183
rect -813 -1225 -811 -1222
rect -916 -1237 -836 -1235
rect -838 -1248 -836 -1237
rect -943 -1260 -939 -1258
rect -919 -1260 -905 -1258
rect -865 -1260 -862 -1258
rect -721 -1229 -719 -1221
rect -82 -1193 -80 -1190
rect -530 -1221 -528 -1217
rect -493 -1221 -491 -1217
rect -377 -1219 -375 -1202
rect -334 -1212 -332 -1198
rect -297 -1212 -295 -1198
rect -185 -1205 -105 -1203
rect -573 -1228 -571 -1224
rect -107 -1216 -105 -1205
rect -212 -1228 -208 -1226
rect -188 -1228 -174 -1226
rect -134 -1228 -131 -1226
rect -334 -1236 -332 -1232
rect -297 -1236 -295 -1232
rect -377 -1243 -375 -1239
rect -107 -1240 -105 -1236
rect -185 -1245 -105 -1243
rect -838 -1272 -836 -1268
rect -916 -1277 -836 -1275
rect -838 -1286 -836 -1277
rect -813 -1279 -811 -1265
rect -721 -1266 -719 -1249
rect -678 -1259 -676 -1245
rect -641 -1259 -639 -1245
rect -107 -1254 -105 -1245
rect -82 -1247 -80 -1233
rect -480 -1258 -478 -1255
rect -443 -1258 -441 -1255
rect -943 -1300 -939 -1298
rect -919 -1300 -905 -1298
rect -865 -1300 -862 -1298
rect -678 -1283 -676 -1279
rect -641 -1283 -639 -1279
rect -523 -1282 -521 -1274
rect -721 -1290 -719 -1286
rect -813 -1303 -811 -1299
rect -212 -1268 -208 -1266
rect -188 -1268 -174 -1266
rect -134 -1268 -131 -1266
rect -82 -1271 -80 -1267
rect -107 -1278 -105 -1274
rect -838 -1310 -836 -1306
rect -523 -1319 -521 -1302
rect -480 -1312 -478 -1298
rect -443 -1312 -441 -1298
rect -480 -1336 -478 -1332
rect -443 -1336 -441 -1332
rect -523 -1343 -521 -1339
rect -840 -1364 -838 -1361
rect -803 -1364 -801 -1361
rect -883 -1388 -881 -1380
rect -679 -1374 -677 -1371
rect -642 -1374 -640 -1371
rect -722 -1398 -720 -1390
rect -883 -1425 -881 -1408
rect -840 -1418 -838 -1404
rect -803 -1418 -801 -1404
rect -722 -1435 -720 -1418
rect -679 -1428 -677 -1414
rect -642 -1428 -640 -1414
rect -840 -1442 -838 -1438
rect -803 -1442 -801 -1438
rect -883 -1449 -881 -1445
rect -679 -1452 -677 -1448
rect -642 -1452 -640 -1448
rect -722 -1459 -720 -1455
rect -776 -1559 -774 -1556
rect -739 -1559 -737 -1556
rect -819 -1583 -817 -1575
rect -615 -1569 -613 -1566
rect -578 -1569 -576 -1566
rect -658 -1593 -656 -1585
rect -819 -1620 -817 -1603
rect -776 -1613 -774 -1599
rect -739 -1613 -737 -1599
rect -658 -1630 -656 -1613
rect -615 -1623 -613 -1609
rect -578 -1623 -576 -1609
rect -776 -1637 -774 -1633
rect -739 -1637 -737 -1633
rect -819 -1644 -817 -1640
rect -615 -1647 -613 -1643
rect -578 -1647 -576 -1643
rect -658 -1654 -656 -1650
rect -775 -1677 -773 -1674
rect -738 -1677 -736 -1674
rect -818 -1701 -816 -1693
rect -818 -1738 -816 -1721
rect -775 -1731 -773 -1717
rect -738 -1731 -736 -1717
rect -775 -1755 -773 -1751
rect -738 -1755 -736 -1751
rect -818 -1762 -816 -1758
rect -937 -1813 -935 -1810
rect -900 -1813 -898 -1810
rect -980 -1837 -978 -1829
rect -980 -1874 -978 -1857
rect -937 -1867 -935 -1853
rect -900 -1867 -898 -1853
rect -937 -1891 -935 -1887
rect -900 -1891 -898 -1887
rect -980 -1898 -978 -1894
rect -592 -1895 -590 -1892
rect -555 -1895 -553 -1892
rect -635 -1919 -633 -1911
rect -875 -1926 -873 -1923
rect -978 -1938 -898 -1936
rect -900 -1949 -898 -1938
rect -1005 -1961 -1001 -1959
rect -981 -1961 -967 -1959
rect -927 -1961 -924 -1959
rect -744 -1927 -742 -1924
rect -707 -1927 -705 -1924
rect -787 -1951 -785 -1943
rect -900 -1973 -898 -1969
rect -978 -1978 -898 -1976
rect -900 -1987 -898 -1978
rect -875 -1980 -873 -1966
rect -417 -1926 -415 -1923
rect -380 -1926 -378 -1923
rect -635 -1956 -633 -1939
rect -592 -1949 -590 -1935
rect -555 -1949 -553 -1935
rect -1005 -2001 -1001 -1999
rect -981 -2001 -967 -1999
rect -927 -2001 -924 -1999
rect -787 -1988 -785 -1971
rect -744 -1981 -742 -1967
rect -707 -1981 -705 -1967
rect -460 -1950 -458 -1942
rect -592 -1973 -590 -1969
rect -555 -1973 -553 -1969
rect -635 -1980 -633 -1976
rect -875 -2004 -873 -2000
rect -900 -2011 -898 -2007
rect -460 -1987 -458 -1970
rect -417 -1980 -415 -1966
rect -380 -1980 -378 -1966
rect -744 -2005 -742 -2001
rect -707 -2005 -705 -2001
rect -417 -2004 -415 -2000
rect -380 -2004 -378 -2000
rect -787 -2012 -785 -2008
rect -460 -2011 -458 -2007
rect -554 -2085 -552 -2082
rect -517 -2085 -515 -2082
rect -597 -2109 -595 -2101
rect -696 -2112 -694 -2109
rect -659 -2112 -657 -2109
rect -739 -2136 -737 -2128
rect -597 -2146 -595 -2129
rect -554 -2139 -552 -2125
rect -517 -2139 -515 -2125
rect -739 -2173 -737 -2156
rect -696 -2166 -694 -2152
rect -659 -2166 -657 -2152
rect -554 -2163 -552 -2159
rect -517 -2163 -515 -2159
rect -597 -2170 -595 -2166
rect -696 -2190 -694 -2186
rect -659 -2190 -657 -2186
rect -739 -2197 -737 -2193
rect -1065 -2219 -1063 -2216
rect -1028 -2219 -1026 -2216
rect -1108 -2243 -1106 -2235
rect -904 -2229 -902 -2226
rect -867 -2229 -865 -2226
rect -947 -2253 -945 -2245
rect -1108 -2280 -1106 -2263
rect -1065 -2273 -1063 -2259
rect -1028 -2273 -1026 -2259
rect -947 -2290 -945 -2273
rect -904 -2283 -902 -2269
rect -867 -2283 -865 -2269
rect -1065 -2297 -1063 -2293
rect -1028 -2297 -1026 -2293
rect -1108 -2304 -1106 -2300
rect -904 -2307 -902 -2303
rect -867 -2307 -865 -2303
rect -947 -2314 -945 -2310
rect -1010 -2351 -1008 -2348
rect -973 -2351 -971 -2348
rect -1053 -2375 -1051 -2367
rect -849 -2361 -847 -2358
rect -812 -2361 -810 -2358
rect -892 -2385 -890 -2377
rect -1053 -2412 -1051 -2395
rect -1010 -2405 -1008 -2391
rect -973 -2405 -971 -2391
rect -892 -2422 -890 -2405
rect -849 -2415 -847 -2401
rect -812 -2415 -810 -2401
rect -1010 -2429 -1008 -2425
rect -973 -2429 -971 -2425
rect -1053 -2436 -1051 -2432
rect -849 -2439 -847 -2435
rect -812 -2439 -810 -2435
rect -892 -2446 -890 -2442
rect -1009 -2469 -1007 -2466
rect -972 -2469 -970 -2466
rect -1052 -2493 -1050 -2485
rect -1052 -2530 -1050 -2513
rect -1009 -2523 -1007 -2509
rect -972 -2523 -970 -2509
rect -1009 -2547 -1007 -2543
rect -972 -2547 -970 -2543
rect -1052 -2554 -1050 -2550
rect -808 -2598 -806 -2595
rect -771 -2598 -769 -2595
rect -851 -2622 -849 -2614
rect -683 -2629 -681 -2626
rect -646 -2629 -644 -2626
rect -851 -2659 -849 -2642
rect -808 -2652 -806 -2638
rect -771 -2652 -769 -2638
rect -726 -2653 -724 -2645
rect -808 -2676 -806 -2672
rect -771 -2676 -769 -2672
rect -851 -2683 -849 -2679
rect -726 -2690 -724 -2673
rect -683 -2683 -681 -2669
rect -646 -2683 -644 -2669
rect -683 -2707 -681 -2703
rect -646 -2707 -644 -2703
rect -726 -2714 -724 -2710
rect -991 -2725 -989 -2722
rect -954 -2725 -952 -2722
rect -1034 -2749 -1032 -2741
rect -830 -2735 -828 -2732
rect -793 -2735 -791 -2732
rect -873 -2759 -871 -2751
rect -1034 -2786 -1032 -2769
rect -991 -2779 -989 -2765
rect -954 -2779 -952 -2765
rect -873 -2796 -871 -2779
rect -830 -2789 -828 -2775
rect -793 -2789 -791 -2775
rect -991 -2803 -989 -2799
rect -954 -2803 -952 -2799
rect -1034 -2810 -1032 -2806
rect -830 -2813 -828 -2809
rect -793 -2813 -791 -2809
rect -873 -2820 -871 -2816
<< polycontact >>
rect -381 -252 -377 -248
rect -381 -269 -377 -265
rect -381 -286 -377 -282
rect -282 -287 -278 -283
rect -381 -309 -377 -305
rect -914 -379 -909 -374
rect -870 -409 -866 -405
rect -833 -409 -829 -405
rect -569 -461 -564 -456
rect -907 -487 -903 -483
rect -907 -504 -903 -500
rect -525 -491 -521 -487
rect -488 -491 -484 -487
rect -907 -521 -903 -517
rect -808 -522 -804 -518
rect -717 -523 -712 -518
rect -907 -544 -903 -540
rect -371 -506 -367 -502
rect -371 -523 -367 -519
rect -371 -540 -367 -536
rect -272 -541 -268 -537
rect -673 -553 -669 -549
rect -636 -553 -632 -549
rect -371 -563 -367 -559
rect -922 -651 -917 -646
rect -878 -681 -874 -677
rect -841 -681 -837 -677
rect -577 -733 -572 -728
rect -381 -748 -376 -743
rect -533 -763 -529 -759
rect -496 -763 -492 -759
rect -725 -795 -720 -790
rect -915 -811 -911 -807
rect -915 -828 -911 -824
rect -337 -778 -333 -774
rect -300 -778 -296 -774
rect -184 -778 -180 -774
rect -184 -795 -180 -791
rect -184 -812 -180 -808
rect -85 -813 -81 -809
rect -681 -825 -677 -821
rect -644 -825 -640 -821
rect -915 -845 -911 -841
rect -816 -846 -812 -842
rect -915 -868 -911 -864
rect -184 -835 -180 -831
rect -725 -911 -720 -906
rect -564 -921 -559 -916
rect -681 -941 -677 -937
rect -644 -941 -640 -937
rect -520 -951 -516 -947
rect -483 -951 -479 -947
rect -923 -1082 -918 -1077
rect -879 -1112 -875 -1108
rect -842 -1112 -838 -1108
rect -578 -1164 -573 -1159
rect -382 -1179 -377 -1174
rect -534 -1194 -530 -1190
rect -497 -1194 -493 -1190
rect -916 -1241 -912 -1237
rect -916 -1258 -912 -1254
rect -726 -1226 -721 -1221
rect -338 -1209 -334 -1205
rect -301 -1209 -297 -1205
rect -185 -1209 -181 -1205
rect -185 -1226 -181 -1222
rect -185 -1243 -181 -1239
rect -86 -1244 -82 -1240
rect -916 -1275 -912 -1271
rect -817 -1276 -813 -1272
rect -682 -1256 -678 -1252
rect -645 -1256 -641 -1252
rect -916 -1298 -912 -1294
rect -528 -1279 -523 -1274
rect -185 -1266 -181 -1262
rect -484 -1309 -480 -1305
rect -447 -1309 -443 -1305
rect -888 -1385 -883 -1380
rect -727 -1395 -722 -1390
rect -844 -1415 -840 -1411
rect -807 -1415 -803 -1411
rect -683 -1425 -679 -1421
rect -646 -1425 -642 -1421
rect -824 -1580 -819 -1575
rect -663 -1590 -658 -1585
rect -780 -1610 -776 -1606
rect -743 -1610 -739 -1606
rect -619 -1620 -615 -1616
rect -582 -1620 -578 -1616
rect -823 -1698 -818 -1693
rect -779 -1728 -775 -1724
rect -742 -1728 -738 -1724
rect -985 -1834 -980 -1829
rect -941 -1864 -937 -1860
rect -904 -1864 -900 -1860
rect -640 -1916 -635 -1911
rect -978 -1942 -974 -1938
rect -978 -1959 -974 -1955
rect -792 -1948 -787 -1943
rect -978 -1976 -974 -1972
rect -879 -1977 -875 -1973
rect -596 -1946 -592 -1942
rect -559 -1946 -555 -1942
rect -465 -1947 -460 -1942
rect -978 -1999 -974 -1995
rect -748 -1978 -744 -1974
rect -711 -1978 -707 -1974
rect -421 -1977 -417 -1973
rect -384 -1977 -380 -1973
rect -602 -2106 -597 -2101
rect -744 -2133 -739 -2128
rect -558 -2136 -554 -2132
rect -521 -2136 -517 -2132
rect -700 -2163 -696 -2159
rect -663 -2163 -659 -2159
rect -1113 -2240 -1108 -2235
rect -952 -2250 -947 -2245
rect -1069 -2270 -1065 -2266
rect -1032 -2270 -1028 -2266
rect -908 -2280 -904 -2276
rect -871 -2280 -867 -2276
rect -1058 -2372 -1053 -2367
rect -897 -2382 -892 -2377
rect -1014 -2402 -1010 -2398
rect -977 -2402 -973 -2398
rect -853 -2412 -849 -2408
rect -816 -2412 -812 -2408
rect -1057 -2490 -1052 -2485
rect -1013 -2520 -1009 -2516
rect -976 -2520 -972 -2516
rect -856 -2619 -851 -2614
rect -812 -2649 -808 -2645
rect -775 -2649 -771 -2645
rect -731 -2650 -726 -2645
rect -687 -2680 -683 -2676
rect -650 -2680 -646 -2676
rect -1039 -2746 -1034 -2741
rect -878 -2756 -873 -2751
rect -995 -2776 -991 -2772
rect -958 -2776 -954 -2772
rect -834 -2786 -830 -2782
rect -797 -2786 -793 -2782
<< metal1 >>
rect -289 -224 -265 -221
rect -289 -228 -286 -224
rect -282 -228 -272 -224
rect -268 -228 -265 -224
rect -289 -230 -265 -228
rect -283 -236 -280 -230
rect -1294 -252 -381 -247
rect -415 -259 -409 -258
rect -415 -263 -414 -259
rect -410 -263 -409 -259
rect -415 -264 -409 -263
rect -415 -267 -404 -264
rect -415 -277 -409 -267
rect -381 -265 -377 -252
rect -324 -261 -315 -258
rect -324 -264 -322 -261
rect -330 -265 -322 -264
rect -318 -265 -315 -261
rect -330 -267 -315 -265
rect -384 -276 -370 -273
rect -324 -275 -315 -267
rect -415 -281 -414 -277
rect -410 -281 -409 -277
rect -415 -282 -409 -281
rect -381 -282 -377 -276
rect -324 -279 -322 -275
rect -318 -279 -315 -275
rect -324 -282 -315 -279
rect -308 -289 -304 -279
rect -1354 -294 -304 -289
rect -299 -283 -296 -279
rect -274 -283 -271 -276
rect -299 -287 -282 -283
rect -274 -287 -263 -283
rect -415 -299 -409 -298
rect -415 -303 -414 -299
rect -410 -303 -409 -299
rect -415 -304 -409 -303
rect -415 -307 -404 -304
rect -415 -317 -409 -307
rect -381 -305 -377 -294
rect -299 -297 -296 -287
rect -274 -290 -271 -287
rect -324 -301 -315 -298
rect -324 -304 -322 -301
rect -330 -305 -322 -304
rect -318 -305 -315 -301
rect -330 -307 -315 -305
rect -384 -316 -370 -313
rect -324 -315 -315 -307
rect -1278 -323 -775 -318
rect -415 -321 -414 -317
rect -410 -321 -409 -317
rect -415 -322 -409 -321
rect -1308 -599 -1289 -594
rect -1278 -917 -1273 -323
rect -877 -346 -853 -343
rect -877 -350 -874 -346
rect -870 -350 -860 -346
rect -856 -350 -853 -346
rect -877 -352 -853 -350
rect -840 -346 -816 -343
rect -840 -350 -837 -346
rect -833 -350 -823 -346
rect -819 -350 -816 -346
rect -840 -352 -816 -350
rect -871 -358 -868 -352
rect -834 -358 -831 -352
rect -961 -379 -951 -374
rect -946 -379 -914 -374
rect -914 -404 -910 -402
rect -971 -409 -960 -404
rect -955 -409 -910 -404
rect -780 -390 -775 -323
rect -381 -333 -377 -316
rect -324 -319 -322 -315
rect -318 -319 -315 -315
rect -324 -322 -315 -319
rect -283 -315 -280 -310
rect -289 -316 -265 -315
rect -308 -333 -304 -317
rect -289 -320 -288 -316
rect -284 -320 -270 -316
rect -266 -320 -265 -316
rect -289 -321 -265 -320
rect -381 -337 -304 -333
rect -906 -405 -902 -402
rect -862 -405 -859 -398
rect -825 -405 -822 -398
rect -906 -409 -870 -405
rect -862 -409 -833 -405
rect -906 -419 -902 -409
rect -862 -412 -859 -409
rect -825 -410 -780 -405
rect -775 -410 -592 -405
rect -825 -412 -822 -410
rect -871 -437 -868 -432
rect -834 -437 -831 -432
rect -877 -438 -853 -437
rect -914 -446 -910 -439
rect -877 -442 -876 -438
rect -872 -442 -858 -438
rect -854 -442 -853 -438
rect -877 -443 -853 -442
rect -840 -438 -816 -437
rect -840 -442 -839 -438
rect -835 -442 -821 -438
rect -817 -442 -816 -438
rect -840 -443 -816 -442
rect -921 -451 -895 -446
rect -598 -456 -592 -410
rect -532 -428 -508 -425
rect -532 -432 -529 -428
rect -525 -432 -515 -428
rect -511 -432 -508 -428
rect -532 -434 -508 -432
rect -495 -428 -471 -425
rect -495 -432 -492 -428
rect -488 -432 -478 -428
rect -474 -432 -471 -428
rect -495 -434 -471 -432
rect -526 -440 -523 -434
rect -489 -440 -486 -434
rect -815 -459 -791 -456
rect -815 -463 -812 -459
rect -808 -463 -798 -459
rect -794 -463 -791 -459
rect -598 -461 -569 -456
rect -815 -465 -791 -463
rect -809 -471 -806 -465
rect -946 -487 -907 -483
rect -941 -494 -935 -493
rect -941 -498 -940 -494
rect -936 -498 -935 -494
rect -941 -499 -935 -498
rect -941 -502 -930 -499
rect -941 -512 -935 -502
rect -907 -500 -903 -487
rect -850 -496 -841 -493
rect -850 -499 -848 -496
rect -856 -500 -848 -499
rect -844 -500 -841 -496
rect -856 -502 -841 -500
rect -910 -511 -896 -508
rect -850 -510 -841 -502
rect -941 -516 -940 -512
rect -936 -516 -935 -512
rect -941 -517 -935 -516
rect -907 -517 -903 -511
rect -850 -514 -848 -510
rect -844 -514 -841 -510
rect -850 -517 -841 -514
rect -569 -486 -565 -484
rect -680 -490 -656 -487
rect -680 -494 -677 -490
rect -673 -494 -663 -490
rect -659 -494 -656 -490
rect -680 -496 -656 -494
rect -643 -490 -619 -487
rect -643 -494 -640 -490
rect -636 -494 -626 -490
rect -622 -494 -619 -490
rect -572 -491 -565 -486
rect -561 -487 -557 -484
rect -517 -487 -514 -480
rect -480 -487 -477 -480
rect -279 -478 -255 -475
rect -279 -482 -276 -478
rect -272 -482 -262 -478
rect -258 -482 -255 -478
rect -279 -484 -255 -482
rect -561 -491 -525 -487
rect -517 -491 -488 -487
rect -643 -496 -619 -494
rect -834 -525 -830 -514
rect -955 -529 -830 -525
rect -825 -518 -822 -514
rect -800 -518 -797 -511
rect -674 -502 -671 -496
rect -637 -502 -634 -496
rect -561 -501 -557 -491
rect -517 -494 -514 -491
rect -480 -492 -405 -487
rect -480 -494 -477 -492
rect -825 -522 -808 -518
rect -941 -534 -935 -533
rect -941 -538 -940 -534
rect -936 -538 -935 -534
rect -941 -539 -935 -538
rect -941 -542 -930 -539
rect -941 -552 -935 -542
rect -907 -540 -903 -529
rect -825 -532 -822 -522
rect -800 -523 -743 -518
rect -738 -523 -717 -518
rect -800 -525 -797 -523
rect -850 -536 -841 -533
rect -850 -539 -848 -536
rect -856 -540 -848 -539
rect -844 -540 -841 -536
rect -856 -542 -841 -540
rect -910 -551 -896 -548
rect -850 -550 -841 -542
rect -941 -556 -940 -552
rect -936 -556 -935 -552
rect -941 -557 -935 -556
rect -907 -568 -903 -551
rect -850 -554 -848 -550
rect -844 -554 -841 -550
rect -850 -557 -841 -554
rect -809 -550 -806 -545
rect -717 -548 -713 -546
rect -815 -551 -791 -550
rect -834 -568 -830 -552
rect -815 -555 -814 -551
rect -810 -555 -796 -551
rect -792 -555 -791 -551
rect -763 -553 -713 -548
rect -409 -502 -405 -492
rect -273 -490 -270 -484
rect -409 -506 -371 -502
rect -405 -513 -399 -512
rect -526 -519 -523 -514
rect -489 -519 -486 -514
rect -405 -517 -404 -513
rect -400 -517 -399 -513
rect -405 -518 -399 -517
rect -532 -520 -508 -519
rect -569 -528 -565 -521
rect -532 -524 -531 -520
rect -527 -524 -513 -520
rect -509 -524 -508 -520
rect -532 -525 -508 -524
rect -495 -520 -471 -519
rect -495 -524 -494 -520
rect -490 -524 -476 -520
rect -472 -524 -471 -520
rect -495 -525 -471 -524
rect -405 -521 -394 -518
rect -709 -549 -705 -546
rect -665 -549 -662 -542
rect -628 -549 -625 -542
rect -593 -533 -565 -528
rect -405 -531 -399 -521
rect -371 -519 -367 -506
rect -314 -515 -305 -512
rect -314 -518 -312 -515
rect -320 -519 -312 -518
rect -308 -519 -305 -515
rect -320 -521 -305 -519
rect -374 -530 -360 -527
rect -314 -529 -305 -521
rect -593 -549 -588 -533
rect -405 -535 -404 -531
rect -400 -535 -399 -531
rect -405 -536 -399 -535
rect -371 -536 -367 -530
rect -314 -533 -312 -529
rect -308 -533 -305 -529
rect -314 -536 -305 -533
rect -298 -543 -294 -533
rect -441 -548 -294 -543
rect -289 -537 -286 -533
rect -264 -537 -261 -530
rect -289 -541 -272 -537
rect -264 -541 -253 -537
rect -709 -553 -673 -549
rect -665 -553 -636 -549
rect -628 -553 -588 -549
rect -405 -553 -399 -552
rect -815 -556 -791 -555
rect -709 -563 -705 -553
rect -665 -556 -662 -553
rect -628 -556 -625 -553
rect -907 -572 -830 -568
rect -405 -557 -404 -553
rect -400 -557 -399 -553
rect -405 -558 -399 -557
rect -405 -561 -394 -558
rect -405 -571 -399 -561
rect -371 -559 -367 -548
rect -289 -551 -286 -541
rect -264 -544 -261 -541
rect -314 -555 -305 -552
rect -314 -558 -312 -555
rect -320 -559 -312 -558
rect -308 -559 -305 -555
rect -320 -561 -305 -559
rect -374 -570 -360 -567
rect -314 -569 -305 -561
rect -405 -575 -404 -571
rect -400 -575 -399 -571
rect -405 -576 -399 -575
rect -674 -581 -671 -576
rect -637 -581 -634 -576
rect -680 -582 -656 -581
rect -717 -590 -713 -583
rect -680 -586 -679 -582
rect -675 -586 -661 -582
rect -657 -586 -656 -582
rect -680 -587 -656 -586
rect -643 -582 -619 -581
rect -643 -586 -642 -582
rect -638 -586 -624 -582
rect -620 -586 -619 -582
rect -643 -587 -619 -586
rect -371 -587 -367 -570
rect -314 -573 -312 -569
rect -308 -573 -305 -569
rect -314 -576 -305 -573
rect -273 -569 -270 -564
rect -279 -570 -255 -569
rect -298 -587 -294 -571
rect -279 -574 -278 -570
rect -274 -574 -260 -570
rect -256 -574 -255 -570
rect -279 -575 -255 -574
rect -724 -595 -698 -590
rect -371 -591 -294 -587
rect -1269 -605 -785 -601
rect -1269 -917 -1264 -605
rect -885 -618 -861 -615
rect -885 -622 -882 -618
rect -878 -622 -868 -618
rect -864 -622 -861 -618
rect -885 -624 -861 -622
rect -848 -618 -824 -615
rect -848 -622 -845 -618
rect -841 -622 -831 -618
rect -827 -622 -824 -618
rect -848 -624 -824 -622
rect -879 -630 -876 -624
rect -842 -630 -839 -624
rect -969 -651 -959 -646
rect -954 -651 -922 -646
rect -922 -676 -918 -674
rect -979 -681 -968 -676
rect -963 -681 -918 -676
rect -914 -677 -910 -674
rect -870 -677 -867 -670
rect -833 -677 -830 -670
rect -794 -677 -787 -605
rect -914 -681 -878 -677
rect -870 -681 -841 -677
rect -833 -681 -600 -677
rect -914 -691 -910 -681
rect -870 -684 -867 -681
rect -833 -684 -830 -681
rect -823 -682 -600 -681
rect -879 -709 -876 -704
rect -842 -709 -839 -704
rect -885 -710 -861 -709
rect -922 -718 -918 -711
rect -885 -714 -884 -710
rect -880 -714 -866 -710
rect -862 -714 -861 -710
rect -885 -715 -861 -714
rect -848 -710 -824 -709
rect -848 -714 -847 -710
rect -843 -714 -829 -710
rect -825 -714 -824 -710
rect -848 -715 -824 -714
rect -929 -723 -903 -718
rect -606 -728 -600 -682
rect -540 -700 -516 -697
rect -540 -704 -537 -700
rect -533 -704 -523 -700
rect -519 -704 -516 -700
rect -540 -706 -516 -704
rect -503 -700 -479 -697
rect -503 -704 -500 -700
rect -496 -704 -486 -700
rect -482 -704 -479 -700
rect -503 -706 -479 -704
rect -534 -712 -531 -706
rect -497 -712 -494 -706
rect -606 -733 -577 -728
rect -577 -758 -573 -756
rect -688 -762 -664 -759
rect -688 -766 -685 -762
rect -681 -766 -671 -762
rect -667 -766 -664 -762
rect -1218 -771 -785 -766
rect -688 -768 -664 -766
rect -651 -762 -627 -759
rect -651 -766 -648 -762
rect -644 -766 -634 -762
rect -630 -766 -627 -762
rect -580 -763 -573 -758
rect -344 -715 -320 -712
rect -344 -719 -341 -715
rect -337 -719 -327 -715
rect -323 -719 -320 -715
rect -344 -721 -320 -719
rect -307 -715 -283 -712
rect -307 -719 -304 -715
rect -300 -719 -290 -715
rect -286 -719 -283 -715
rect -307 -721 -283 -719
rect -338 -727 -335 -721
rect -301 -727 -298 -721
rect -569 -759 -565 -756
rect -525 -759 -522 -752
rect -488 -759 -485 -752
rect -411 -748 -381 -743
rect -411 -759 -406 -748
rect -569 -763 -533 -759
rect -525 -763 -496 -759
rect -488 -763 -406 -759
rect -651 -768 -627 -766
rect -823 -783 -799 -780
rect -823 -787 -820 -783
rect -816 -787 -806 -783
rect -802 -787 -799 -783
rect -823 -789 -799 -787
rect -817 -795 -814 -789
rect -790 -790 -785 -771
rect -682 -774 -679 -768
rect -645 -774 -642 -768
rect -569 -773 -565 -763
rect -525 -766 -522 -763
rect -488 -766 -485 -763
rect -790 -795 -725 -790
rect -954 -811 -915 -807
rect -949 -818 -943 -817
rect -949 -822 -948 -818
rect -944 -822 -943 -818
rect -949 -823 -943 -822
rect -949 -826 -938 -823
rect -949 -836 -943 -826
rect -915 -824 -911 -811
rect -858 -820 -849 -817
rect -858 -823 -856 -820
rect -864 -824 -856 -823
rect -852 -824 -849 -820
rect -864 -826 -849 -824
rect -918 -835 -904 -832
rect -858 -834 -849 -826
rect -949 -840 -948 -836
rect -944 -840 -943 -836
rect -949 -841 -943 -840
rect -915 -841 -911 -835
rect -858 -838 -856 -834
rect -852 -838 -849 -834
rect -858 -841 -849 -838
rect -725 -820 -721 -818
rect -842 -849 -838 -838
rect -963 -853 -838 -849
rect -833 -842 -830 -838
rect -808 -842 -805 -835
rect -780 -825 -771 -820
rect -766 -825 -721 -820
rect -381 -773 -377 -771
rect -384 -778 -377 -773
rect -92 -750 -68 -747
rect -92 -754 -89 -750
rect -85 -754 -75 -750
rect -71 -754 -68 -750
rect -92 -756 -68 -754
rect -373 -774 -369 -771
rect -329 -774 -326 -767
rect -292 -774 -289 -767
rect -86 -762 -83 -756
rect -373 -778 -337 -774
rect -329 -778 -300 -774
rect -292 -778 -184 -774
rect -534 -791 -531 -786
rect -497 -791 -494 -786
rect -373 -788 -369 -778
rect -329 -781 -326 -778
rect -292 -781 -289 -778
rect -540 -792 -516 -791
rect -577 -800 -573 -793
rect -540 -796 -539 -792
rect -535 -796 -521 -792
rect -517 -796 -516 -792
rect -540 -797 -516 -796
rect -503 -792 -479 -791
rect -503 -796 -502 -792
rect -498 -796 -484 -792
rect -480 -796 -479 -792
rect -503 -797 -479 -796
rect -717 -821 -713 -818
rect -673 -821 -670 -814
rect -636 -821 -633 -814
rect -601 -805 -573 -800
rect -601 -821 -596 -805
rect -218 -785 -212 -784
rect -218 -789 -217 -785
rect -213 -789 -212 -785
rect -218 -790 -212 -789
rect -218 -793 -207 -790
rect -338 -806 -335 -801
rect -301 -806 -298 -801
rect -218 -803 -212 -793
rect -184 -791 -180 -778
rect -127 -787 -118 -784
rect -127 -790 -125 -787
rect -133 -791 -125 -790
rect -121 -791 -118 -787
rect -133 -793 -118 -791
rect -187 -802 -173 -799
rect -127 -801 -118 -793
rect -344 -807 -320 -806
rect -381 -815 -377 -808
rect -344 -811 -343 -807
rect -339 -811 -325 -807
rect -321 -811 -320 -807
rect -344 -812 -320 -811
rect -307 -807 -283 -806
rect -307 -811 -306 -807
rect -302 -811 -288 -807
rect -284 -811 -283 -807
rect -218 -807 -217 -803
rect -213 -807 -212 -803
rect -218 -808 -212 -807
rect -184 -808 -180 -802
rect -127 -805 -125 -801
rect -121 -805 -118 -801
rect -127 -808 -118 -805
rect -307 -812 -283 -811
rect -111 -815 -107 -805
rect -717 -825 -681 -821
rect -673 -825 -644 -821
rect -636 -825 -596 -821
rect -474 -820 -377 -815
rect -233 -820 -107 -815
rect -102 -809 -99 -805
rect -77 -809 -74 -802
rect -102 -813 -85 -809
rect -77 -813 -66 -809
rect -780 -842 -775 -825
rect -717 -835 -713 -825
rect -673 -828 -670 -825
rect -636 -828 -633 -825
rect -833 -846 -816 -842
rect -949 -858 -943 -857
rect -949 -862 -948 -858
rect -944 -862 -943 -858
rect -949 -863 -943 -862
rect -949 -866 -938 -863
rect -949 -876 -943 -866
rect -915 -864 -911 -853
rect -833 -856 -830 -846
rect -808 -847 -775 -842
rect -808 -849 -805 -847
rect -858 -860 -849 -857
rect -858 -863 -856 -860
rect -864 -864 -856 -863
rect -852 -864 -849 -860
rect -864 -866 -849 -864
rect -918 -875 -904 -872
rect -858 -874 -849 -866
rect -949 -880 -948 -876
rect -944 -880 -943 -876
rect -949 -881 -943 -880
rect -915 -892 -911 -875
rect -858 -878 -856 -874
rect -852 -878 -849 -874
rect -858 -881 -849 -878
rect -682 -853 -679 -848
rect -645 -853 -642 -848
rect -688 -854 -664 -853
rect -725 -862 -721 -855
rect -688 -858 -687 -854
rect -683 -858 -669 -854
rect -665 -858 -664 -854
rect -688 -859 -664 -858
rect -651 -854 -627 -853
rect -651 -858 -650 -854
rect -646 -858 -632 -854
rect -628 -858 -627 -854
rect -651 -859 -627 -858
rect -732 -867 -706 -862
rect -817 -874 -814 -869
rect -474 -870 -468 -820
rect -218 -825 -212 -824
rect -218 -829 -217 -825
rect -213 -829 -212 -825
rect -218 -830 -212 -829
rect -218 -833 -207 -830
rect -218 -843 -212 -833
rect -184 -831 -180 -820
rect -102 -823 -99 -813
rect -77 -816 -74 -813
rect -127 -827 -118 -824
rect -127 -830 -125 -827
rect -133 -831 -125 -830
rect -121 -831 -118 -827
rect -133 -833 -118 -831
rect -187 -842 -173 -839
rect -127 -841 -118 -833
rect -218 -847 -217 -843
rect -213 -847 -212 -843
rect -218 -848 -212 -847
rect -184 -859 -180 -842
rect -127 -845 -125 -841
rect -121 -845 -118 -841
rect -127 -848 -118 -845
rect -86 -841 -83 -836
rect -92 -842 -68 -841
rect -111 -859 -107 -843
rect -92 -846 -91 -842
rect -87 -846 -73 -842
rect -69 -846 -68 -842
rect -92 -847 -68 -846
rect -184 -863 -107 -859
rect -474 -874 -428 -870
rect -823 -875 -799 -874
rect -842 -892 -838 -876
rect -823 -879 -822 -875
rect -818 -879 -804 -875
rect -800 -879 -799 -875
rect -823 -880 -799 -879
rect -688 -878 -664 -875
rect -688 -882 -685 -878
rect -681 -882 -671 -878
rect -667 -882 -664 -878
rect -688 -884 -664 -882
rect -651 -878 -627 -875
rect -651 -882 -648 -878
rect -644 -882 -634 -878
rect -630 -882 -627 -878
rect -651 -884 -627 -882
rect -915 -896 -838 -892
rect -682 -890 -679 -884
rect -645 -890 -642 -884
rect -527 -888 -503 -885
rect -804 -911 -725 -906
rect -804 -927 -799 -911
rect -1354 -932 -799 -927
rect -725 -936 -721 -934
rect -1294 -941 -721 -936
rect -527 -892 -524 -888
rect -520 -892 -510 -888
rect -506 -892 -503 -888
rect -527 -894 -503 -892
rect -490 -888 -466 -885
rect -490 -892 -487 -888
rect -483 -892 -473 -888
rect -469 -892 -466 -888
rect -490 -894 -466 -892
rect -521 -900 -518 -894
rect -484 -900 -481 -894
rect -717 -937 -713 -934
rect -673 -937 -670 -930
rect -636 -937 -633 -930
rect -593 -921 -564 -916
rect -593 -937 -587 -921
rect -717 -941 -681 -937
rect -673 -941 -644 -937
rect -636 -941 -587 -937
rect -1278 -1565 -1273 -953
rect -717 -951 -713 -941
rect -673 -944 -670 -941
rect -636 -944 -633 -941
rect -1269 -1565 -1264 -953
rect -564 -946 -560 -944
rect -587 -951 -560 -946
rect -556 -947 -552 -944
rect -512 -947 -509 -940
rect -475 -947 -472 -940
rect -432 -947 -428 -874
rect -556 -951 -520 -947
rect -512 -951 -483 -947
rect -475 -951 -428 -947
rect -682 -969 -679 -964
rect -645 -969 -642 -964
rect -688 -970 -664 -969
rect -725 -978 -721 -971
rect -688 -974 -687 -970
rect -683 -974 -669 -970
rect -665 -974 -664 -970
rect -688 -975 -664 -974
rect -651 -970 -627 -969
rect -651 -974 -650 -970
rect -646 -974 -632 -970
rect -628 -974 -627 -970
rect -651 -975 -627 -974
rect -732 -983 -706 -978
rect -587 -987 -582 -951
rect -556 -961 -552 -951
rect -512 -954 -509 -951
rect -475 -954 -472 -951
rect -1255 -992 -582 -987
rect -521 -979 -518 -974
rect -484 -979 -481 -974
rect -527 -980 -503 -979
rect -564 -988 -560 -981
rect -527 -984 -526 -980
rect -522 -984 -508 -980
rect -504 -984 -503 -980
rect -527 -985 -503 -984
rect -490 -980 -466 -979
rect -490 -984 -489 -980
rect -485 -984 -471 -980
rect -467 -984 -466 -980
rect -490 -985 -466 -984
rect -571 -993 -545 -988
rect -886 -1049 -862 -1046
rect -886 -1053 -883 -1049
rect -879 -1053 -869 -1049
rect -865 -1053 -862 -1049
rect -886 -1055 -862 -1053
rect -849 -1049 -825 -1046
rect -849 -1053 -846 -1049
rect -842 -1053 -832 -1049
rect -828 -1053 -825 -1049
rect -849 -1055 -825 -1053
rect -880 -1061 -877 -1055
rect -843 -1061 -840 -1055
rect -970 -1082 -960 -1077
rect -955 -1082 -923 -1077
rect -923 -1107 -919 -1105
rect -980 -1112 -969 -1107
rect -964 -1112 -919 -1107
rect -915 -1108 -911 -1105
rect -871 -1108 -868 -1101
rect -834 -1108 -831 -1101
rect -915 -1112 -879 -1108
rect -871 -1112 -842 -1108
rect -915 -1122 -911 -1112
rect -871 -1115 -868 -1112
rect -834 -1113 -601 -1108
rect -834 -1115 -831 -1113
rect -880 -1140 -877 -1135
rect -843 -1140 -840 -1135
rect -886 -1141 -862 -1140
rect -923 -1149 -919 -1142
rect -886 -1145 -885 -1141
rect -881 -1145 -867 -1141
rect -863 -1145 -862 -1141
rect -886 -1146 -862 -1145
rect -849 -1141 -825 -1140
rect -849 -1145 -848 -1141
rect -844 -1145 -830 -1141
rect -826 -1145 -825 -1141
rect -849 -1146 -825 -1145
rect -930 -1154 -904 -1149
rect -607 -1159 -601 -1113
rect -541 -1131 -517 -1128
rect -541 -1135 -538 -1131
rect -534 -1135 -524 -1131
rect -520 -1135 -517 -1131
rect -541 -1137 -517 -1135
rect -504 -1131 -480 -1128
rect -504 -1135 -501 -1131
rect -497 -1135 -487 -1131
rect -483 -1135 -480 -1131
rect -504 -1137 -480 -1135
rect -535 -1143 -532 -1137
rect -498 -1143 -495 -1137
rect -607 -1164 -578 -1159
rect -1251 -1187 -784 -1182
rect -824 -1213 -800 -1210
rect -824 -1217 -821 -1213
rect -817 -1217 -807 -1213
rect -803 -1217 -800 -1213
rect -824 -1219 -800 -1217
rect -818 -1225 -815 -1219
rect -789 -1221 -784 -1187
rect -578 -1189 -574 -1187
rect -689 -1193 -665 -1190
rect -689 -1197 -686 -1193
rect -682 -1197 -672 -1193
rect -668 -1197 -665 -1193
rect -689 -1199 -665 -1197
rect -652 -1193 -628 -1190
rect -652 -1197 -649 -1193
rect -645 -1197 -635 -1193
rect -631 -1197 -628 -1193
rect -581 -1194 -574 -1189
rect -345 -1146 -321 -1143
rect -345 -1150 -342 -1146
rect -338 -1150 -328 -1146
rect -324 -1150 -321 -1146
rect -345 -1152 -321 -1150
rect -308 -1146 -284 -1143
rect -308 -1150 -305 -1146
rect -301 -1150 -291 -1146
rect -287 -1150 -284 -1146
rect -308 -1152 -284 -1150
rect -339 -1158 -336 -1152
rect -302 -1158 -299 -1152
rect -570 -1190 -566 -1187
rect -526 -1190 -523 -1183
rect -489 -1190 -486 -1183
rect -412 -1179 -382 -1174
rect -412 -1190 -407 -1179
rect -570 -1194 -534 -1190
rect -526 -1194 -497 -1190
rect -489 -1194 -407 -1190
rect -652 -1199 -628 -1197
rect -683 -1205 -680 -1199
rect -646 -1205 -643 -1199
rect -570 -1204 -566 -1194
rect -526 -1197 -523 -1194
rect -489 -1197 -486 -1194
rect -955 -1241 -916 -1237
rect -950 -1248 -944 -1247
rect -950 -1252 -949 -1248
rect -945 -1252 -944 -1248
rect -950 -1253 -944 -1252
rect -950 -1256 -939 -1253
rect -950 -1266 -944 -1256
rect -916 -1254 -912 -1241
rect -859 -1250 -850 -1247
rect -859 -1253 -857 -1250
rect -865 -1254 -857 -1253
rect -853 -1254 -850 -1250
rect -865 -1256 -850 -1254
rect -919 -1265 -905 -1262
rect -859 -1264 -850 -1256
rect -950 -1270 -949 -1266
rect -945 -1270 -944 -1266
rect -950 -1271 -944 -1270
rect -916 -1271 -912 -1265
rect -859 -1268 -857 -1264
rect -853 -1268 -850 -1264
rect -859 -1271 -850 -1268
rect -789 -1226 -726 -1221
rect -726 -1251 -722 -1249
rect -843 -1279 -839 -1268
rect -964 -1283 -839 -1279
rect -834 -1272 -831 -1268
rect -809 -1272 -806 -1265
rect -791 -1256 -772 -1251
rect -767 -1256 -722 -1251
rect -382 -1204 -378 -1202
rect -385 -1209 -378 -1204
rect -93 -1181 -69 -1178
rect -93 -1185 -90 -1181
rect -86 -1185 -76 -1181
rect -72 -1185 -69 -1181
rect -93 -1187 -69 -1185
rect -374 -1205 -370 -1202
rect -330 -1205 -327 -1198
rect -293 -1205 -290 -1198
rect -87 -1193 -84 -1187
rect -374 -1209 -338 -1205
rect -330 -1209 -301 -1205
rect -293 -1209 -185 -1205
rect -535 -1222 -532 -1217
rect -498 -1222 -495 -1217
rect -374 -1219 -370 -1209
rect -330 -1212 -327 -1209
rect -293 -1212 -290 -1209
rect -541 -1223 -517 -1222
rect -578 -1231 -574 -1224
rect -541 -1227 -540 -1223
rect -536 -1227 -522 -1223
rect -518 -1227 -517 -1223
rect -541 -1228 -517 -1227
rect -504 -1223 -480 -1222
rect -504 -1227 -503 -1223
rect -499 -1227 -485 -1223
rect -481 -1227 -480 -1223
rect -504 -1228 -480 -1227
rect -718 -1252 -714 -1249
rect -674 -1252 -671 -1245
rect -637 -1252 -634 -1245
rect -602 -1236 -574 -1231
rect -602 -1252 -597 -1236
rect -219 -1216 -213 -1215
rect -219 -1220 -218 -1216
rect -214 -1220 -213 -1216
rect -219 -1221 -213 -1220
rect -219 -1224 -208 -1221
rect -339 -1237 -336 -1232
rect -302 -1237 -299 -1232
rect -219 -1234 -213 -1224
rect -185 -1222 -181 -1209
rect -128 -1218 -119 -1215
rect -128 -1221 -126 -1218
rect -134 -1222 -126 -1221
rect -122 -1222 -119 -1218
rect -134 -1224 -119 -1222
rect -188 -1233 -174 -1230
rect -128 -1232 -119 -1224
rect -345 -1238 -321 -1237
rect -491 -1246 -467 -1243
rect -491 -1250 -488 -1246
rect -484 -1250 -474 -1246
rect -470 -1250 -467 -1246
rect -491 -1252 -467 -1250
rect -454 -1246 -430 -1243
rect -382 -1246 -378 -1239
rect -345 -1242 -344 -1238
rect -340 -1242 -326 -1238
rect -322 -1242 -321 -1238
rect -345 -1243 -321 -1242
rect -308 -1238 -284 -1237
rect -308 -1242 -307 -1238
rect -303 -1242 -289 -1238
rect -285 -1242 -284 -1238
rect -219 -1238 -218 -1234
rect -214 -1238 -213 -1234
rect -219 -1239 -213 -1238
rect -185 -1239 -181 -1233
rect -128 -1236 -126 -1232
rect -122 -1236 -119 -1232
rect -128 -1239 -119 -1236
rect -308 -1243 -284 -1242
rect -112 -1246 -108 -1236
rect -454 -1250 -451 -1246
rect -447 -1250 -437 -1246
rect -433 -1250 -430 -1246
rect -454 -1252 -430 -1250
rect -422 -1251 -378 -1246
rect -214 -1251 -108 -1246
rect -103 -1240 -100 -1236
rect -78 -1240 -75 -1233
rect -103 -1244 -86 -1240
rect -78 -1244 -67 -1240
rect -718 -1256 -682 -1252
rect -674 -1256 -645 -1252
rect -637 -1256 -597 -1252
rect -791 -1272 -786 -1256
rect -718 -1266 -714 -1256
rect -674 -1259 -671 -1256
rect -637 -1259 -634 -1256
rect -834 -1276 -817 -1272
rect -950 -1288 -944 -1287
rect -950 -1292 -949 -1288
rect -945 -1292 -944 -1288
rect -950 -1293 -944 -1292
rect -950 -1296 -939 -1293
rect -950 -1306 -944 -1296
rect -916 -1294 -912 -1283
rect -834 -1286 -831 -1276
rect -809 -1277 -786 -1272
rect -809 -1279 -806 -1277
rect -859 -1290 -850 -1287
rect -859 -1293 -857 -1290
rect -865 -1294 -857 -1293
rect -853 -1294 -850 -1290
rect -865 -1296 -850 -1294
rect -919 -1305 -905 -1302
rect -859 -1304 -850 -1296
rect -950 -1310 -949 -1306
rect -945 -1310 -944 -1306
rect -950 -1311 -944 -1310
rect -916 -1322 -912 -1305
rect -859 -1308 -857 -1304
rect -853 -1308 -850 -1304
rect -859 -1311 -850 -1308
rect -485 -1258 -482 -1252
rect -448 -1258 -445 -1252
rect -595 -1279 -528 -1274
rect -683 -1284 -680 -1279
rect -646 -1284 -643 -1279
rect -689 -1285 -665 -1284
rect -726 -1293 -722 -1286
rect -689 -1289 -688 -1285
rect -684 -1289 -670 -1285
rect -666 -1289 -665 -1285
rect -689 -1290 -665 -1289
rect -652 -1285 -628 -1284
rect -652 -1289 -651 -1285
rect -647 -1289 -633 -1285
rect -629 -1289 -628 -1285
rect -652 -1290 -628 -1289
rect -733 -1298 -707 -1293
rect -818 -1304 -815 -1299
rect -824 -1305 -800 -1304
rect -843 -1322 -839 -1306
rect -824 -1309 -823 -1305
rect -819 -1309 -805 -1305
rect -801 -1309 -800 -1305
rect -824 -1310 -800 -1309
rect -916 -1326 -839 -1322
rect -851 -1352 -827 -1349
rect -851 -1356 -848 -1352
rect -844 -1356 -834 -1352
rect -830 -1356 -827 -1352
rect -851 -1358 -827 -1356
rect -814 -1352 -790 -1349
rect -814 -1356 -811 -1352
rect -807 -1356 -797 -1352
rect -793 -1356 -790 -1352
rect -814 -1358 -790 -1356
rect -845 -1364 -842 -1358
rect -808 -1364 -805 -1358
rect -690 -1362 -666 -1359
rect -1224 -1385 -888 -1380
rect -888 -1410 -884 -1408
rect -1255 -1415 -884 -1410
rect -690 -1366 -687 -1362
rect -683 -1366 -673 -1362
rect -669 -1366 -666 -1362
rect -690 -1368 -666 -1366
rect -653 -1362 -629 -1359
rect -653 -1366 -650 -1362
rect -646 -1366 -636 -1362
rect -632 -1366 -629 -1362
rect -653 -1368 -629 -1366
rect -684 -1374 -681 -1368
rect -647 -1374 -644 -1368
rect -880 -1411 -876 -1408
rect -836 -1411 -833 -1404
rect -799 -1411 -796 -1404
rect -756 -1395 -727 -1390
rect -756 -1411 -750 -1395
rect -880 -1415 -844 -1411
rect -836 -1415 -807 -1411
rect -799 -1415 -750 -1411
rect -880 -1425 -876 -1415
rect -836 -1418 -833 -1415
rect -799 -1418 -796 -1415
rect -727 -1420 -723 -1418
rect -750 -1425 -723 -1420
rect -719 -1421 -715 -1418
rect -675 -1421 -672 -1414
rect -638 -1421 -635 -1414
rect -595 -1421 -591 -1279
rect -528 -1304 -524 -1302
rect -531 -1309 -524 -1304
rect -520 -1305 -516 -1302
rect -476 -1305 -473 -1298
rect -439 -1305 -436 -1298
rect -422 -1305 -417 -1251
rect -219 -1256 -213 -1255
rect -219 -1260 -218 -1256
rect -214 -1260 -213 -1256
rect -219 -1261 -213 -1260
rect -219 -1264 -208 -1261
rect -219 -1274 -213 -1264
rect -185 -1262 -181 -1251
rect -103 -1254 -100 -1244
rect -78 -1247 -75 -1244
rect -128 -1258 -119 -1255
rect -128 -1261 -126 -1258
rect -134 -1262 -126 -1261
rect -122 -1262 -119 -1258
rect -134 -1264 -119 -1262
rect -188 -1273 -174 -1270
rect -128 -1272 -119 -1264
rect -219 -1278 -218 -1274
rect -214 -1278 -213 -1274
rect -219 -1279 -213 -1278
rect -185 -1290 -181 -1273
rect -128 -1276 -126 -1272
rect -122 -1276 -119 -1272
rect -128 -1279 -119 -1276
rect -87 -1272 -84 -1267
rect -93 -1273 -69 -1272
rect -112 -1290 -108 -1274
rect -93 -1277 -92 -1273
rect -88 -1277 -74 -1273
rect -70 -1277 -69 -1273
rect -93 -1278 -69 -1277
rect -185 -1294 -108 -1290
rect -520 -1309 -484 -1305
rect -476 -1309 -447 -1305
rect -439 -1309 -417 -1305
rect -520 -1319 -516 -1309
rect -476 -1312 -473 -1309
rect -439 -1312 -436 -1309
rect -429 -1310 -417 -1309
rect -485 -1337 -482 -1332
rect -448 -1337 -445 -1332
rect -491 -1338 -467 -1337
rect -528 -1346 -524 -1339
rect -491 -1342 -490 -1338
rect -486 -1342 -472 -1338
rect -468 -1342 -467 -1338
rect -491 -1343 -467 -1342
rect -454 -1338 -430 -1337
rect -454 -1342 -453 -1338
rect -449 -1342 -435 -1338
rect -431 -1342 -430 -1338
rect -454 -1343 -430 -1342
rect -719 -1425 -683 -1421
rect -675 -1425 -646 -1421
rect -638 -1425 -591 -1421
rect -543 -1351 -524 -1346
rect -845 -1443 -842 -1438
rect -808 -1443 -805 -1438
rect -851 -1444 -827 -1443
rect -888 -1452 -884 -1445
rect -851 -1448 -850 -1444
rect -846 -1448 -832 -1444
rect -828 -1448 -827 -1444
rect -851 -1449 -827 -1448
rect -814 -1444 -790 -1443
rect -814 -1448 -813 -1444
rect -809 -1448 -795 -1444
rect -791 -1448 -790 -1444
rect -814 -1449 -790 -1448
rect -895 -1457 -869 -1452
rect -750 -1471 -745 -1425
rect -719 -1435 -715 -1425
rect -675 -1428 -672 -1425
rect -638 -1428 -635 -1425
rect -684 -1453 -681 -1448
rect -647 -1453 -644 -1448
rect -690 -1454 -666 -1453
rect -727 -1462 -723 -1455
rect -690 -1458 -689 -1454
rect -685 -1458 -671 -1454
rect -667 -1458 -666 -1454
rect -690 -1459 -666 -1458
rect -653 -1454 -629 -1453
rect -653 -1458 -652 -1454
rect -648 -1458 -634 -1454
rect -630 -1458 -629 -1454
rect -653 -1459 -629 -1458
rect -734 -1467 -708 -1462
rect -1248 -1476 -745 -1471
rect -543 -1544 -536 -1351
rect -787 -1547 -763 -1544
rect -787 -1551 -784 -1547
rect -780 -1551 -770 -1547
rect -766 -1551 -763 -1547
rect -787 -1553 -763 -1551
rect -750 -1547 -726 -1544
rect -750 -1551 -747 -1547
rect -743 -1551 -733 -1547
rect -729 -1551 -726 -1547
rect -750 -1553 -726 -1551
rect -781 -1559 -778 -1553
rect -744 -1559 -741 -1553
rect -626 -1557 -602 -1554
rect -1354 -1580 -824 -1575
rect -824 -1605 -820 -1603
rect -1294 -1610 -820 -1605
rect -626 -1561 -623 -1557
rect -619 -1561 -609 -1557
rect -605 -1561 -602 -1557
rect -626 -1563 -602 -1561
rect -589 -1557 -565 -1554
rect -589 -1561 -586 -1557
rect -582 -1561 -572 -1557
rect -568 -1561 -565 -1557
rect -589 -1563 -565 -1561
rect -620 -1569 -617 -1563
rect -583 -1569 -580 -1563
rect -816 -1606 -812 -1603
rect -772 -1606 -769 -1599
rect -735 -1606 -732 -1599
rect -692 -1590 -663 -1585
rect -692 -1606 -686 -1590
rect -816 -1610 -780 -1606
rect -772 -1610 -743 -1606
rect -735 -1610 -686 -1606
rect -1278 -2515 -1273 -1619
rect -1269 -2318 -1264 -1619
rect -816 -1620 -812 -1610
rect -772 -1613 -769 -1610
rect -735 -1613 -732 -1610
rect -663 -1615 -659 -1613
rect -693 -1620 -659 -1615
rect -655 -1616 -651 -1613
rect -611 -1616 -608 -1609
rect -574 -1616 -571 -1609
rect -543 -1616 -537 -1544
rect -655 -1620 -619 -1616
rect -611 -1620 -582 -1616
rect -574 -1620 -537 -1616
rect -781 -1638 -778 -1633
rect -744 -1638 -741 -1633
rect -787 -1639 -763 -1638
rect -824 -1647 -820 -1640
rect -787 -1643 -786 -1639
rect -782 -1643 -768 -1639
rect -764 -1643 -763 -1639
rect -787 -1644 -763 -1643
rect -750 -1639 -726 -1638
rect -750 -1643 -749 -1639
rect -745 -1643 -731 -1639
rect -727 -1643 -726 -1639
rect -750 -1644 -726 -1643
rect -831 -1652 -805 -1647
rect -786 -1665 -762 -1662
rect -786 -1669 -783 -1665
rect -779 -1669 -769 -1665
rect -765 -1669 -762 -1665
rect -786 -1671 -762 -1669
rect -749 -1665 -725 -1662
rect -749 -1669 -746 -1665
rect -742 -1669 -732 -1665
rect -728 -1669 -725 -1665
rect -749 -1671 -725 -1669
rect -780 -1677 -777 -1671
rect -743 -1677 -740 -1671
rect -1255 -1698 -823 -1693
rect -823 -1723 -819 -1721
rect -1224 -1728 -819 -1723
rect -815 -1724 -811 -1721
rect -771 -1724 -768 -1717
rect -734 -1724 -731 -1717
rect -693 -1724 -686 -1620
rect -655 -1630 -651 -1620
rect -611 -1623 -608 -1620
rect -574 -1623 -571 -1620
rect -620 -1648 -617 -1643
rect -583 -1648 -580 -1643
rect -626 -1649 -602 -1648
rect -663 -1657 -659 -1650
rect -626 -1653 -625 -1649
rect -621 -1653 -607 -1649
rect -603 -1653 -602 -1649
rect -626 -1654 -602 -1653
rect -589 -1649 -565 -1648
rect -589 -1653 -588 -1649
rect -584 -1653 -570 -1649
rect -566 -1653 -565 -1649
rect -589 -1654 -565 -1653
rect -670 -1662 -644 -1657
rect -815 -1728 -779 -1724
rect -771 -1728 -742 -1724
rect -734 -1728 -686 -1724
rect -815 -1738 -811 -1728
rect -771 -1731 -768 -1728
rect -734 -1731 -731 -1728
rect -780 -1756 -777 -1751
rect -743 -1756 -740 -1751
rect -786 -1757 -762 -1756
rect -823 -1765 -819 -1758
rect -786 -1761 -785 -1757
rect -781 -1761 -767 -1757
rect -763 -1761 -762 -1757
rect -786 -1762 -762 -1761
rect -749 -1757 -725 -1756
rect -749 -1761 -748 -1757
rect -744 -1761 -730 -1757
rect -726 -1761 -725 -1757
rect -749 -1762 -725 -1761
rect -830 -1770 -804 -1765
rect -948 -1801 -924 -1798
rect -948 -1805 -945 -1801
rect -941 -1805 -931 -1801
rect -927 -1805 -924 -1801
rect -948 -1807 -924 -1805
rect -911 -1801 -887 -1798
rect -911 -1805 -908 -1801
rect -904 -1805 -894 -1801
rect -890 -1805 -887 -1801
rect -911 -1807 -887 -1805
rect -942 -1813 -939 -1807
rect -905 -1813 -902 -1807
rect -1032 -1834 -1022 -1829
rect -1017 -1834 -985 -1829
rect -985 -1859 -981 -1857
rect -1042 -1864 -1031 -1859
rect -1026 -1864 -981 -1859
rect -977 -1860 -973 -1857
rect -933 -1860 -930 -1853
rect -896 -1860 -893 -1853
rect -977 -1864 -941 -1860
rect -933 -1864 -904 -1860
rect -977 -1874 -973 -1864
rect -933 -1867 -930 -1864
rect -896 -1865 -663 -1860
rect -896 -1867 -893 -1865
rect -942 -1892 -939 -1887
rect -905 -1892 -902 -1887
rect -948 -1893 -924 -1892
rect -985 -1901 -981 -1894
rect -948 -1897 -947 -1893
rect -943 -1897 -929 -1893
rect -925 -1897 -924 -1893
rect -948 -1898 -924 -1897
rect -911 -1893 -887 -1892
rect -911 -1897 -910 -1893
rect -906 -1897 -892 -1893
rect -888 -1897 -887 -1893
rect -911 -1898 -887 -1897
rect -992 -1906 -966 -1901
rect -669 -1911 -663 -1865
rect -603 -1883 -579 -1880
rect -603 -1887 -600 -1883
rect -596 -1887 -586 -1883
rect -582 -1887 -579 -1883
rect -603 -1889 -579 -1887
rect -566 -1883 -542 -1880
rect -566 -1887 -563 -1883
rect -559 -1887 -549 -1883
rect -545 -1887 -542 -1883
rect -566 -1889 -542 -1887
rect -597 -1895 -594 -1889
rect -560 -1895 -557 -1889
rect -886 -1914 -862 -1911
rect -886 -1918 -883 -1914
rect -879 -1918 -869 -1914
rect -865 -1918 -862 -1914
rect -886 -1920 -862 -1918
rect -755 -1915 -731 -1912
rect -755 -1919 -752 -1915
rect -748 -1919 -738 -1915
rect -734 -1919 -731 -1915
rect -880 -1926 -877 -1920
rect -755 -1921 -731 -1919
rect -718 -1915 -694 -1912
rect -718 -1919 -715 -1915
rect -711 -1919 -701 -1915
rect -697 -1919 -694 -1915
rect -669 -1916 -640 -1911
rect -718 -1921 -694 -1919
rect -1017 -1942 -978 -1938
rect -1012 -1949 -1006 -1948
rect -1012 -1953 -1011 -1949
rect -1007 -1953 -1006 -1949
rect -1012 -1954 -1006 -1953
rect -1012 -1957 -1001 -1954
rect -1012 -1967 -1006 -1957
rect -978 -1955 -974 -1942
rect -921 -1951 -912 -1948
rect -921 -1954 -919 -1951
rect -927 -1955 -919 -1954
rect -915 -1955 -912 -1951
rect -927 -1957 -912 -1955
rect -981 -1966 -967 -1963
rect -921 -1965 -912 -1957
rect -1012 -1971 -1011 -1967
rect -1007 -1971 -1006 -1967
rect -1012 -1972 -1006 -1971
rect -978 -1972 -974 -1966
rect -921 -1969 -919 -1965
rect -915 -1969 -912 -1965
rect -921 -1972 -912 -1969
rect -749 -1927 -746 -1921
rect -712 -1927 -709 -1921
rect -827 -1948 -792 -1943
rect -905 -1980 -901 -1969
rect -1026 -1984 -901 -1980
rect -896 -1973 -893 -1969
rect -871 -1973 -868 -1966
rect -792 -1973 -788 -1971
rect -896 -1977 -879 -1973
rect -1012 -1989 -1006 -1988
rect -1012 -1993 -1011 -1989
rect -1007 -1993 -1006 -1989
rect -1012 -1994 -1006 -1993
rect -1012 -1997 -1001 -1994
rect -1012 -2007 -1006 -1997
rect -978 -1995 -974 -1984
rect -896 -1987 -893 -1977
rect -871 -1978 -847 -1973
rect -842 -1978 -788 -1973
rect -640 -1941 -636 -1939
rect -643 -1946 -636 -1941
rect -428 -1914 -404 -1911
rect -428 -1918 -425 -1914
rect -421 -1918 -411 -1914
rect -407 -1918 -404 -1914
rect -428 -1920 -404 -1918
rect -391 -1914 -367 -1911
rect -391 -1918 -388 -1914
rect -384 -1918 -374 -1914
rect -370 -1918 -367 -1914
rect -391 -1920 -367 -1918
rect -632 -1942 -628 -1939
rect -588 -1942 -585 -1935
rect -551 -1942 -548 -1935
rect -422 -1926 -419 -1920
rect -385 -1926 -382 -1920
rect -632 -1946 -596 -1942
rect -588 -1946 -559 -1942
rect -632 -1956 -628 -1946
rect -588 -1949 -585 -1946
rect -551 -1947 -465 -1942
rect -551 -1949 -548 -1947
rect -784 -1974 -780 -1971
rect -740 -1974 -737 -1967
rect -703 -1974 -700 -1967
rect -784 -1978 -748 -1974
rect -740 -1978 -711 -1974
rect -703 -1978 -669 -1974
rect -871 -1980 -868 -1978
rect -921 -1991 -912 -1988
rect -921 -1994 -919 -1991
rect -927 -1995 -919 -1994
rect -915 -1995 -912 -1991
rect -927 -1997 -912 -1995
rect -981 -2006 -967 -2003
rect -921 -2005 -912 -1997
rect -1012 -2011 -1011 -2007
rect -1007 -2011 -1006 -2007
rect -1012 -2012 -1006 -2011
rect -978 -2023 -974 -2006
rect -921 -2009 -919 -2005
rect -915 -2009 -912 -2005
rect -921 -2012 -912 -2009
rect -784 -1988 -780 -1978
rect -740 -1981 -737 -1978
rect -703 -1981 -700 -1978
rect -880 -2005 -877 -2000
rect -886 -2006 -862 -2005
rect -905 -2023 -901 -2007
rect -886 -2010 -885 -2006
rect -881 -2010 -867 -2006
rect -863 -2010 -862 -2006
rect -886 -2011 -862 -2010
rect -674 -1983 -669 -1978
rect -597 -1974 -594 -1969
rect -560 -1974 -557 -1969
rect -465 -1972 -461 -1970
rect -603 -1975 -579 -1974
rect -640 -1983 -636 -1976
rect -603 -1979 -602 -1975
rect -598 -1979 -584 -1975
rect -580 -1979 -579 -1975
rect -603 -1980 -579 -1979
rect -566 -1975 -542 -1974
rect -566 -1979 -565 -1975
rect -561 -1979 -547 -1975
rect -543 -1979 -542 -1975
rect -468 -1977 -461 -1972
rect -457 -1973 -453 -1970
rect -413 -1973 -410 -1966
rect -376 -1973 -373 -1966
rect -457 -1977 -421 -1973
rect -413 -1977 -384 -1973
rect -376 -1977 -358 -1973
rect -566 -1980 -542 -1979
rect -674 -1988 -636 -1983
rect -457 -1987 -453 -1977
rect -413 -1980 -410 -1977
rect -376 -1980 -373 -1977
rect -749 -2006 -746 -2001
rect -712 -2006 -709 -2001
rect -755 -2007 -731 -2006
rect -792 -2015 -788 -2008
rect -755 -2011 -754 -2007
rect -750 -2011 -736 -2007
rect -732 -2011 -731 -2007
rect -755 -2012 -731 -2011
rect -718 -2007 -694 -2006
rect -718 -2011 -717 -2007
rect -713 -2011 -699 -2007
rect -695 -2011 -694 -2007
rect -718 -2012 -694 -2011
rect -422 -2005 -419 -2000
rect -385 -2005 -382 -2000
rect -428 -2006 -404 -2005
rect -465 -2014 -461 -2007
rect -428 -2010 -427 -2006
rect -423 -2010 -409 -2006
rect -405 -2010 -404 -2006
rect -428 -2011 -404 -2010
rect -391 -2006 -367 -2005
rect -391 -2010 -390 -2006
rect -386 -2010 -372 -2006
rect -368 -2010 -367 -2006
rect -391 -2011 -367 -2010
rect -799 -2020 -773 -2015
rect -978 -2027 -901 -2023
rect -494 -2021 -461 -2014
rect -565 -2073 -541 -2070
rect -565 -2077 -562 -2073
rect -558 -2077 -548 -2073
rect -544 -2077 -541 -2073
rect -565 -2079 -541 -2077
rect -528 -2073 -504 -2070
rect -528 -2077 -525 -2073
rect -521 -2077 -511 -2073
rect -507 -2077 -504 -2073
rect -528 -2079 -504 -2077
rect -559 -2085 -556 -2079
rect -522 -2085 -519 -2079
rect -707 -2100 -683 -2097
rect -707 -2104 -704 -2100
rect -700 -2104 -690 -2100
rect -686 -2104 -683 -2100
rect -707 -2106 -683 -2104
rect -670 -2100 -646 -2097
rect -670 -2104 -667 -2100
rect -663 -2104 -653 -2100
rect -649 -2104 -646 -2100
rect -670 -2106 -646 -2104
rect -638 -2106 -602 -2101
rect -701 -2112 -698 -2106
rect -664 -2112 -661 -2106
rect -821 -2133 -744 -2128
rect -821 -2187 -816 -2133
rect -744 -2158 -740 -2156
rect -747 -2163 -740 -2158
rect -736 -2159 -732 -2156
rect -692 -2159 -689 -2152
rect -655 -2159 -652 -2152
rect -638 -2159 -633 -2106
rect -602 -2131 -598 -2129
rect -605 -2136 -598 -2131
rect -594 -2132 -590 -2129
rect -550 -2132 -547 -2125
rect -513 -2132 -510 -2125
rect -494 -2132 -486 -2021
rect -594 -2136 -558 -2132
rect -550 -2136 -521 -2132
rect -513 -2136 -486 -2132
rect -594 -2146 -590 -2136
rect -550 -2139 -547 -2136
rect -513 -2139 -510 -2136
rect -736 -2163 -700 -2159
rect -692 -2163 -663 -2159
rect -655 -2163 -633 -2159
rect -736 -2173 -732 -2163
rect -692 -2166 -689 -2163
rect -655 -2166 -652 -2163
rect -645 -2164 -633 -2163
rect -1076 -2207 -1052 -2204
rect -1076 -2211 -1073 -2207
rect -1069 -2211 -1059 -2207
rect -1055 -2211 -1052 -2207
rect -1076 -2213 -1052 -2211
rect -1039 -2207 -1015 -2204
rect -1039 -2211 -1036 -2207
rect -1032 -2211 -1022 -2207
rect -1018 -2211 -1015 -2207
rect -1039 -2213 -1015 -2211
rect -1070 -2219 -1067 -2213
rect -1033 -2219 -1030 -2213
rect -915 -2217 -891 -2214
rect -1179 -2240 -1113 -2235
rect -1113 -2265 -1109 -2263
rect -1224 -2270 -1109 -2265
rect -915 -2221 -912 -2217
rect -908 -2221 -898 -2217
rect -894 -2221 -891 -2217
rect -915 -2223 -891 -2221
rect -878 -2217 -854 -2214
rect -878 -2221 -875 -2217
rect -871 -2221 -861 -2217
rect -857 -2221 -854 -2217
rect -878 -2223 -854 -2221
rect -909 -2229 -906 -2223
rect -872 -2229 -869 -2223
rect -1105 -2266 -1101 -2263
rect -1061 -2266 -1058 -2259
rect -1024 -2266 -1021 -2259
rect -981 -2250 -952 -2245
rect -981 -2266 -975 -2250
rect -1105 -2270 -1069 -2266
rect -1061 -2270 -1032 -2266
rect -1024 -2270 -975 -2266
rect -1105 -2280 -1101 -2270
rect -1061 -2273 -1058 -2270
rect -1024 -2273 -1021 -2270
rect -952 -2275 -948 -2273
rect -975 -2280 -948 -2275
rect -944 -2276 -940 -2273
rect -900 -2276 -897 -2269
rect -863 -2276 -860 -2269
rect -822 -2276 -816 -2187
rect -559 -2164 -556 -2159
rect -522 -2164 -519 -2159
rect -565 -2165 -541 -2164
rect -602 -2173 -598 -2166
rect -565 -2169 -564 -2165
rect -560 -2169 -546 -2165
rect -542 -2169 -541 -2165
rect -565 -2170 -541 -2169
rect -528 -2165 -504 -2164
rect -528 -2169 -527 -2165
rect -523 -2169 -509 -2165
rect -505 -2169 -504 -2165
rect -528 -2170 -504 -2169
rect -628 -2178 -598 -2173
rect -701 -2191 -698 -2186
rect -664 -2191 -661 -2186
rect -707 -2192 -683 -2191
rect -744 -2200 -740 -2193
rect -707 -2196 -706 -2192
rect -702 -2196 -688 -2192
rect -684 -2196 -683 -2192
rect -707 -2197 -683 -2196
rect -670 -2192 -646 -2191
rect -670 -2196 -669 -2192
rect -665 -2196 -651 -2192
rect -647 -2196 -646 -2192
rect -670 -2197 -646 -2196
rect -768 -2205 -740 -2200
rect -768 -2210 -761 -2205
rect -944 -2280 -908 -2276
rect -900 -2280 -871 -2276
rect -863 -2280 -816 -2276
rect -777 -2215 -761 -2210
rect -1070 -2298 -1067 -2293
rect -1033 -2298 -1030 -2293
rect -1076 -2299 -1052 -2298
rect -1113 -2307 -1109 -2300
rect -1076 -2303 -1075 -2299
rect -1071 -2303 -1057 -2299
rect -1053 -2303 -1052 -2299
rect -1076 -2304 -1052 -2303
rect -1039 -2299 -1015 -2298
rect -1039 -2303 -1038 -2299
rect -1034 -2303 -1020 -2299
rect -1016 -2303 -1015 -2299
rect -1039 -2304 -1015 -2303
rect -1120 -2312 -1094 -2307
rect -975 -2318 -970 -2280
rect -944 -2290 -940 -2280
rect -900 -2283 -897 -2280
rect -863 -2283 -860 -2280
rect -909 -2308 -906 -2303
rect -872 -2308 -869 -2303
rect -915 -2309 -891 -2308
rect -952 -2317 -948 -2310
rect -915 -2313 -914 -2309
rect -910 -2313 -896 -2309
rect -892 -2313 -891 -2309
rect -915 -2314 -891 -2313
rect -878 -2309 -854 -2308
rect -878 -2313 -877 -2309
rect -873 -2313 -859 -2309
rect -855 -2313 -854 -2309
rect -878 -2314 -854 -2313
rect -1269 -2323 -970 -2318
rect -959 -2322 -933 -2317
rect -1021 -2339 -997 -2336
rect -1021 -2343 -1018 -2339
rect -1014 -2343 -1004 -2339
rect -1000 -2343 -997 -2339
rect -1021 -2345 -997 -2343
rect -984 -2339 -960 -2336
rect -984 -2343 -981 -2339
rect -977 -2343 -967 -2339
rect -963 -2343 -960 -2339
rect -984 -2345 -960 -2343
rect -1015 -2351 -1012 -2345
rect -978 -2351 -975 -2345
rect -860 -2349 -836 -2346
rect -1179 -2372 -1058 -2367
rect -1058 -2397 -1054 -2395
rect -1224 -2402 -1054 -2397
rect -860 -2353 -857 -2349
rect -853 -2353 -843 -2349
rect -839 -2353 -836 -2349
rect -860 -2355 -836 -2353
rect -823 -2349 -799 -2346
rect -823 -2353 -820 -2349
rect -816 -2353 -806 -2349
rect -802 -2353 -799 -2349
rect -823 -2355 -799 -2353
rect -854 -2361 -851 -2355
rect -817 -2361 -814 -2355
rect -1050 -2398 -1046 -2395
rect -1006 -2398 -1003 -2391
rect -969 -2398 -966 -2391
rect -926 -2382 -897 -2377
rect -926 -2398 -920 -2382
rect -1050 -2402 -1014 -2398
rect -1006 -2402 -977 -2398
rect -969 -2402 -920 -2398
rect -1050 -2412 -1046 -2402
rect -1006 -2405 -1003 -2402
rect -969 -2405 -966 -2402
rect -897 -2407 -893 -2405
rect -927 -2412 -893 -2407
rect -889 -2408 -885 -2405
rect -845 -2408 -842 -2401
rect -808 -2408 -805 -2401
rect -777 -2408 -770 -2215
rect -889 -2412 -853 -2408
rect -845 -2412 -816 -2408
rect -808 -2412 -770 -2408
rect -1015 -2430 -1012 -2425
rect -978 -2430 -975 -2425
rect -1021 -2431 -997 -2430
rect -1058 -2439 -1054 -2432
rect -1021 -2435 -1020 -2431
rect -1016 -2435 -1002 -2431
rect -998 -2435 -997 -2431
rect -1021 -2436 -997 -2435
rect -984 -2431 -960 -2430
rect -984 -2435 -983 -2431
rect -979 -2435 -965 -2431
rect -961 -2435 -960 -2431
rect -984 -2436 -960 -2435
rect -1065 -2444 -1039 -2439
rect -1020 -2457 -996 -2454
rect -1020 -2461 -1017 -2457
rect -1013 -2461 -1003 -2457
rect -999 -2461 -996 -2457
rect -1020 -2463 -996 -2461
rect -983 -2457 -959 -2454
rect -983 -2461 -980 -2457
rect -976 -2461 -966 -2457
rect -962 -2461 -959 -2457
rect -983 -2463 -959 -2461
rect -1014 -2469 -1011 -2463
rect -977 -2469 -974 -2463
rect -1255 -2489 -1057 -2485
rect -1260 -2490 -1057 -2489
rect -1057 -2515 -1053 -2513
rect -1278 -2520 -1053 -2515
rect -1049 -2516 -1045 -2513
rect -1005 -2516 -1002 -2509
rect -968 -2516 -965 -2509
rect -927 -2516 -920 -2412
rect -889 -2422 -885 -2412
rect -845 -2415 -842 -2412
rect -808 -2415 -805 -2412
rect -854 -2440 -851 -2435
rect -817 -2440 -814 -2435
rect -860 -2441 -836 -2440
rect -897 -2449 -893 -2442
rect -860 -2445 -859 -2441
rect -855 -2445 -841 -2441
rect -837 -2445 -836 -2441
rect -860 -2446 -836 -2445
rect -823 -2441 -799 -2440
rect -823 -2445 -822 -2441
rect -818 -2445 -804 -2441
rect -800 -2445 -799 -2441
rect -823 -2446 -799 -2445
rect -904 -2454 -878 -2449
rect -1049 -2520 -1013 -2516
rect -1005 -2520 -976 -2516
rect -968 -2520 -920 -2516
rect -1049 -2530 -1045 -2520
rect -1005 -2523 -1002 -2520
rect -968 -2523 -965 -2520
rect -1014 -2548 -1011 -2543
rect -977 -2548 -974 -2543
rect -1020 -2549 -996 -2548
rect -1057 -2557 -1053 -2550
rect -1020 -2553 -1019 -2549
rect -1015 -2553 -1001 -2549
rect -997 -2553 -996 -2549
rect -1020 -2554 -996 -2553
rect -983 -2549 -959 -2548
rect -983 -2553 -982 -2549
rect -978 -2553 -964 -2549
rect -960 -2553 -959 -2549
rect -983 -2554 -959 -2553
rect -1064 -2562 -1038 -2557
rect -819 -2586 -795 -2583
rect -819 -2590 -816 -2586
rect -812 -2590 -802 -2586
rect -798 -2590 -795 -2586
rect -819 -2592 -795 -2590
rect -782 -2586 -758 -2583
rect -782 -2590 -779 -2586
rect -775 -2590 -765 -2586
rect -761 -2590 -758 -2586
rect -782 -2592 -758 -2590
rect -813 -2598 -810 -2592
rect -776 -2598 -773 -2592
rect -1354 -2619 -856 -2614
rect -856 -2644 -852 -2642
rect -1294 -2649 -852 -2644
rect -764 -2608 -758 -2604
rect -694 -2617 -670 -2614
rect -694 -2621 -691 -2617
rect -687 -2621 -677 -2617
rect -673 -2621 -670 -2617
rect -694 -2623 -670 -2621
rect -657 -2617 -633 -2614
rect -657 -2621 -654 -2617
rect -650 -2621 -640 -2617
rect -636 -2621 -633 -2617
rect -657 -2623 -633 -2621
rect -848 -2645 -844 -2642
rect -804 -2645 -801 -2638
rect -767 -2645 -764 -2638
rect -688 -2629 -685 -2623
rect -651 -2629 -648 -2623
rect -848 -2649 -812 -2645
rect -804 -2649 -775 -2645
rect -848 -2659 -844 -2649
rect -804 -2652 -801 -2649
rect -767 -2650 -731 -2645
rect -767 -2652 -764 -2650
rect -813 -2677 -810 -2672
rect -776 -2677 -773 -2672
rect -731 -2675 -727 -2673
rect -819 -2678 -795 -2677
rect -856 -2686 -852 -2679
rect -819 -2682 -818 -2678
rect -814 -2682 -800 -2678
rect -796 -2682 -795 -2678
rect -819 -2683 -795 -2682
rect -782 -2678 -758 -2677
rect -782 -2682 -781 -2678
rect -777 -2682 -763 -2678
rect -759 -2682 -758 -2678
rect -782 -2683 -758 -2682
rect -748 -2680 -727 -2675
rect -723 -2676 -719 -2673
rect -679 -2676 -676 -2669
rect -642 -2676 -639 -2669
rect -628 -2676 -621 -2178
rect -723 -2680 -687 -2676
rect -679 -2680 -650 -2676
rect -642 -2680 -621 -2676
rect -863 -2691 -837 -2686
rect -1002 -2713 -978 -2710
rect -1002 -2717 -999 -2713
rect -995 -2717 -985 -2713
rect -981 -2717 -978 -2713
rect -1002 -2719 -978 -2717
rect -965 -2713 -941 -2710
rect -965 -2717 -962 -2713
rect -958 -2717 -948 -2713
rect -944 -2717 -941 -2713
rect -965 -2719 -941 -2717
rect -996 -2725 -993 -2719
rect -959 -2725 -956 -2719
rect -841 -2723 -817 -2720
rect -1255 -2746 -1039 -2741
rect -1039 -2771 -1035 -2769
rect -1224 -2776 -1035 -2771
rect -841 -2727 -838 -2723
rect -834 -2727 -824 -2723
rect -820 -2727 -817 -2723
rect -841 -2729 -817 -2727
rect -804 -2723 -780 -2720
rect -804 -2727 -801 -2723
rect -797 -2727 -787 -2723
rect -783 -2727 -780 -2723
rect -804 -2729 -780 -2727
rect -835 -2735 -832 -2729
rect -798 -2735 -795 -2729
rect -1031 -2772 -1027 -2769
rect -987 -2772 -984 -2765
rect -950 -2772 -947 -2765
rect -907 -2756 -878 -2751
rect -907 -2772 -901 -2756
rect -1031 -2776 -995 -2772
rect -987 -2776 -958 -2772
rect -950 -2776 -901 -2772
rect -1031 -2786 -1027 -2776
rect -987 -2779 -984 -2776
rect -950 -2779 -947 -2776
rect -878 -2781 -874 -2779
rect -926 -2786 -874 -2781
rect -870 -2782 -866 -2779
rect -826 -2782 -823 -2775
rect -789 -2782 -786 -2775
rect -748 -2782 -742 -2680
rect -723 -2690 -719 -2680
rect -679 -2683 -676 -2680
rect -642 -2683 -639 -2680
rect -688 -2708 -685 -2703
rect -651 -2708 -648 -2703
rect -694 -2709 -670 -2708
rect -731 -2717 -727 -2710
rect -694 -2713 -693 -2709
rect -689 -2713 -675 -2709
rect -671 -2713 -670 -2709
rect -694 -2714 -670 -2713
rect -657 -2709 -633 -2708
rect -657 -2713 -656 -2709
rect -652 -2713 -638 -2709
rect -634 -2713 -633 -2709
rect -657 -2714 -633 -2713
rect -738 -2722 -712 -2717
rect -870 -2786 -834 -2782
rect -826 -2786 -797 -2782
rect -789 -2786 -742 -2782
rect -996 -2804 -993 -2799
rect -959 -2804 -956 -2799
rect -1002 -2805 -978 -2804
rect -1039 -2813 -1035 -2806
rect -1002 -2809 -1001 -2805
rect -997 -2809 -983 -2805
rect -979 -2809 -978 -2805
rect -1002 -2810 -978 -2809
rect -965 -2805 -941 -2804
rect -965 -2809 -964 -2805
rect -960 -2809 -946 -2805
rect -942 -2809 -941 -2805
rect -965 -2810 -941 -2809
rect -1046 -2818 -1020 -2813
rect -926 -2834 -920 -2786
rect -870 -2796 -866 -2786
rect -826 -2789 -823 -2786
rect -789 -2789 -786 -2786
rect -835 -2814 -832 -2809
rect -798 -2814 -795 -2809
rect -841 -2815 -817 -2814
rect -878 -2823 -874 -2816
rect -841 -2819 -840 -2815
rect -836 -2819 -822 -2815
rect -818 -2819 -817 -2815
rect -841 -2820 -817 -2819
rect -804 -2815 -780 -2814
rect -804 -2819 -803 -2815
rect -799 -2819 -785 -2815
rect -781 -2819 -780 -2815
rect -804 -2820 -780 -2819
rect -885 -2828 -859 -2823
rect -1179 -2839 -920 -2834
<< m2contact >>
rect -1299 -252 -1294 -247
rect -1359 -294 -1354 -289
rect -1313 -599 -1308 -594
rect -1289 -599 -1284 -594
rect -951 -379 -946 -374
rect -960 -409 -955 -404
rect -780 -395 -775 -390
rect -780 -410 -775 -405
rect -951 -487 -946 -482
rect -960 -529 -955 -524
rect -743 -523 -738 -518
rect -768 -553 -763 -548
rect -446 -548 -441 -543
rect -1278 -922 -1273 -917
rect -959 -651 -954 -646
rect -968 -681 -963 -676
rect -1223 -771 -1218 -766
rect -959 -811 -954 -806
rect -968 -853 -963 -848
rect -771 -825 -766 -820
rect -238 -820 -233 -815
rect -1269 -922 -1264 -917
rect -1359 -932 -1354 -927
rect -1299 -941 -1294 -936
rect -1278 -953 -1273 -948
rect -1278 -1570 -1273 -1565
rect -1269 -953 -1264 -948
rect -1260 -992 -1255 -987
rect -960 -1082 -955 -1077
rect -969 -1112 -964 -1107
rect -960 -1241 -955 -1236
rect -969 -1283 -964 -1278
rect -772 -1256 -767 -1251
rect -219 -1251 -214 -1246
rect -1229 -1385 -1224 -1380
rect -1260 -1415 -1255 -1410
rect -1269 -1570 -1264 -1565
rect -1359 -1580 -1354 -1575
rect -1299 -1610 -1294 -1605
rect -1278 -1619 -1273 -1614
rect -1269 -1619 -1264 -1614
rect -1260 -1698 -1255 -1693
rect -1229 -1728 -1224 -1723
rect -1022 -1834 -1017 -1829
rect -1031 -1864 -1026 -1859
rect -1022 -1942 -1017 -1937
rect -1031 -1984 -1026 -1979
rect -847 -1978 -842 -1973
rect -1184 -2240 -1179 -2235
rect -1229 -2270 -1224 -2265
rect -1184 -2372 -1179 -2367
rect -1229 -2402 -1224 -2397
rect -1260 -2489 -1255 -2484
rect -1359 -2619 -1354 -2614
rect -1299 -2649 -1294 -2644
rect -1260 -2746 -1255 -2741
rect -1229 -2776 -1224 -2771
rect -1184 -2839 -1179 -2834
<< metal2 >>
rect -1359 -594 -1354 -294
rect -1299 -576 -1294 -252
rect -960 -524 -955 -409
rect -951 -482 -946 -379
rect -780 -405 -775 -395
rect -768 -576 -763 -553
rect -1299 -581 -763 -576
rect -1359 -599 -1313 -594
rect -1359 -927 -1354 -599
rect -1359 -1575 -1354 -932
rect -1359 -2614 -1354 -1580
rect -1299 -766 -1294 -581
rect -743 -594 -738 -523
rect -1284 -599 -738 -594
rect -446 -605 -441 -548
rect -771 -610 -441 -605
rect -1299 -771 -1223 -766
rect -1299 -936 -1294 -771
rect -968 -848 -963 -681
rect -959 -806 -954 -651
rect -771 -820 -766 -610
rect -771 -887 -766 -825
rect -818 -892 -766 -887
rect -818 -911 -812 -892
rect -1260 -916 -812 -911
rect -1299 -1605 -1294 -941
rect -1278 -948 -1273 -922
rect -1269 -948 -1264 -922
rect -1260 -987 -1255 -916
rect -1260 -1410 -1255 -992
rect -238 -1006 -233 -820
rect -772 -1011 -233 -1006
rect -969 -1278 -964 -1112
rect -960 -1236 -955 -1082
rect -772 -1251 -767 -1011
rect -1299 -2644 -1294 -1610
rect -1278 -1614 -1273 -1570
rect -1269 -1614 -1264 -1570
rect -1260 -1693 -1255 -1415
rect -1229 -1301 -1043 -1296
rect -1229 -1380 -1224 -1301
rect -1048 -1330 -1043 -1301
rect -772 -1330 -767 -1256
rect -1048 -1335 -767 -1330
rect -233 -1251 -219 -1246
rect -1260 -2484 -1255 -1698
rect -1260 -2741 -1255 -2489
rect -1229 -1723 -1224 -1385
rect -1229 -2265 -1224 -1728
rect -233 -1782 -228 -1251
rect -847 -1787 -228 -1782
rect -1031 -1979 -1026 -1864
rect -1022 -1937 -1017 -1834
rect -847 -1973 -842 -1787
rect -847 -2048 -842 -1978
rect -1229 -2397 -1224 -2270
rect -1229 -2771 -1224 -2402
rect -1184 -2053 -842 -2048
rect -1184 -2235 -1179 -2053
rect -1184 -2367 -1179 -2240
rect -1184 -2834 -1179 -2372
<< m3contact >>
rect -1269 -1187 -1264 -1182
rect -1251 -1187 -1246 -1182
rect -812 -1113 -807 -1108
rect -1278 -1476 -1273 -1471
rect -1248 -1476 -1243 -1471
rect -827 -1948 -822 -1943
<< metal3 >>
rect -1079 -1028 -807 -1023
rect -1264 -1187 -1251 -1182
rect -1273 -1476 -1248 -1471
rect -1079 -1754 -1074 -1028
rect -812 -1108 -807 -1028
rect -1079 -1759 -864 -1754
rect -869 -1810 -864 -1759
rect -869 -1815 -822 -1810
rect -827 -1943 -822 -1815
<< labels >>
rlabel metal1 -858 -439 -858 -439 8 gnd
rlabel metal1 -863 -351 -863 -351 5 vdd
rlabel metal1 -821 -439 -821 -439 8 gnd
rlabel metal1 -826 -351 -826 -351 5 vdd
rlabel metal1 -911 -449 -911 -449 1 gnd
rlabel metal1 -796 -552 -796 -552 8 gnd
rlabel metal1 -801 -464 -801 -464 5 vdd
rlabel metal1 -937 -512 -937 -512 2 gnd
rlabel metal1 -849 -507 -849 -507 7 vdd
rlabel metal1 -849 -547 -849 -547 7 vdd
rlabel metal1 -937 -552 -937 -552 2 gnd
rlabel metal1 -661 -583 -661 -583 8 gnd
rlabel metal1 -666 -495 -666 -495 5 vdd
rlabel metal1 -624 -583 -624 -583 8 gnd
rlabel metal1 -629 -495 -629 -495 5 vdd
rlabel metal1 -714 -593 -714 -593 1 gnd
rlabel metal1 -569 -489 -569 -489 1 vdd
rlabel metal1 -481 -433 -481 -433 5 vdd
rlabel metal1 -476 -521 -476 -521 8 gnd
rlabel metal1 -518 -433 -518 -433 5 vdd
rlabel metal1 -513 -521 -513 -521 8 gnd
rlabel metal1 -401 -571 -401 -571 2 gnd
rlabel metal1 -313 -566 -313 -566 7 vdd
rlabel metal1 -313 -526 -313 -526 7 vdd
rlabel metal1 -401 -531 -401 -531 2 gnd
rlabel metal1 -265 -483 -265 -483 5 vdd
rlabel metal1 -260 -571 -260 -571 8 gnd
rlabel metal1 -866 -711 -866 -711 8 gnd
rlabel metal1 -871 -623 -871 -623 5 vdd
rlabel metal1 -829 -711 -829 -711 8 gnd
rlabel metal1 -834 -623 -834 -623 5 vdd
rlabel metal1 -919 -721 -919 -721 1 gnd
rlabel metal1 -669 -855 -669 -855 8 gnd
rlabel metal1 -674 -767 -674 -767 5 vdd
rlabel metal1 -632 -855 -632 -855 8 gnd
rlabel metal1 -637 -767 -637 -767 5 vdd
rlabel metal1 -722 -865 -722 -865 1 gnd
rlabel metal1 -577 -761 -577 -761 1 vdd
rlabel metal1 -489 -705 -489 -705 5 vdd
rlabel metal1 -484 -793 -484 -793 8 gnd
rlabel metal1 -526 -705 -526 -705 5 vdd
rlabel metal1 -521 -793 -521 -793 8 gnd
rlabel metal1 -325 -808 -325 -808 8 gnd
rlabel metal1 -330 -720 -330 -720 5 vdd
rlabel metal1 -288 -808 -288 -808 8 gnd
rlabel metal1 -293 -720 -293 -720 5 vdd
rlabel metal1 -381 -776 -381 -776 1 vdd
rlabel metal1 -73 -843 -73 -843 8 gnd
rlabel metal1 -78 -755 -78 -755 5 vdd
rlabel metal1 -214 -803 -214 -803 2 gnd
rlabel metal1 -126 -798 -126 -798 7 vdd
rlabel metal1 -126 -838 -126 -838 7 vdd
rlabel metal1 -214 -843 -214 -843 2 gnd
rlabel metal1 -508 -981 -508 -981 8 gnd
rlabel metal1 -513 -893 -513 -893 5 vdd
rlabel metal1 -471 -981 -471 -981 8 gnd
rlabel metal1 -476 -893 -476 -893 5 vdd
rlabel metal1 -561 -991 -561 -991 1 gnd
rlabel metal1 -722 -981 -722 -981 1 gnd
rlabel metal1 -637 -883 -637 -883 5 vdd
rlabel metal1 -632 -971 -632 -971 8 gnd
rlabel metal1 -674 -883 -674 -883 5 vdd
rlabel metal1 -669 -971 -669 -971 8 gnd
rlabel metal1 -804 -876 -804 -876 8 gnd
rlabel metal1 -809 -788 -809 -788 5 vdd
rlabel metal1 -945 -836 -945 -836 2 gnd
rlabel metal1 -857 -831 -857 -831 7 vdd
rlabel metal1 -857 -871 -857 -871 7 vdd
rlabel metal1 -945 -876 -945 -876 2 gnd
rlabel metal1 -805 -1306 -805 -1306 8 gnd
rlabel metal1 -810 -1218 -810 -1218 5 vdd
rlabel metal1 -946 -1266 -946 -1266 2 gnd
rlabel metal1 -858 -1261 -858 -1261 7 vdd
rlabel metal1 -858 -1301 -858 -1301 7 vdd
rlabel metal1 -946 -1306 -946 -1306 2 gnd
rlabel metal1 -528 -1307 -528 -1307 1 vdd
rlabel metal1 -440 -1251 -440 -1251 5 vdd
rlabel metal1 -435 -1339 -435 -1339 8 gnd
rlabel metal1 -477 -1251 -477 -1251 5 vdd
rlabel metal1 -472 -1339 -472 -1339 8 gnd
rlabel metal1 -215 -1274 -215 -1274 2 gnd
rlabel metal1 -127 -1269 -127 -1269 7 vdd
rlabel metal1 -127 -1229 -127 -1229 7 vdd
rlabel metal1 -215 -1234 -215 -1234 2 gnd
rlabel metal1 -79 -1186 -79 -1186 5 vdd
rlabel metal1 -74 -1274 -74 -1274 8 gnd
rlabel metal1 -382 -1207 -382 -1207 1 vdd
rlabel metal1 -294 -1151 -294 -1151 5 vdd
rlabel metal1 -289 -1239 -289 -1239 8 gnd
rlabel metal1 -331 -1151 -331 -1151 5 vdd
rlabel metal1 -326 -1239 -326 -1239 8 gnd
rlabel metal1 -522 -1224 -522 -1224 8 gnd
rlabel metal1 -527 -1136 -527 -1136 5 vdd
rlabel metal1 -485 -1224 -485 -1224 8 gnd
rlabel metal1 -490 -1136 -490 -1136 5 vdd
rlabel metal1 -578 -1192 -578 -1192 1 vdd
rlabel metal1 -723 -1296 -723 -1296 1 gnd
rlabel metal1 -638 -1198 -638 -1198 5 vdd
rlabel metal1 -633 -1286 -633 -1286 8 gnd
rlabel metal1 -675 -1198 -675 -1198 5 vdd
rlabel metal1 -670 -1286 -670 -1286 8 gnd
rlabel metal1 -920 -1152 -920 -1152 1 gnd
rlabel metal1 -835 -1054 -835 -1054 5 vdd
rlabel metal1 -830 -1142 -830 -1142 8 gnd
rlabel metal1 -872 -1054 -872 -1054 5 vdd
rlabel metal1 -867 -1142 -867 -1142 8 gnd
rlabel metal1 -411 -317 -411 -317 2 gnd
rlabel metal1 -323 -312 -323 -312 7 vdd
rlabel metal1 -323 -272 -323 -272 7 vdd
rlabel metal1 -411 -277 -411 -277 2 gnd
rlabel metal1 -275 -229 -275 -229 5 vdd
rlabel metal1 -270 -317 -270 -317 8 gnd
rlabel metal1 -832 -1445 -832 -1445 8 gnd
rlabel metal1 -837 -1357 -837 -1357 5 vdd
rlabel metal1 -795 -1445 -795 -1445 8 gnd
rlabel metal1 -800 -1357 -800 -1357 5 vdd
rlabel metal1 -885 -1455 -885 -1455 1 gnd
rlabel metal1 -724 -1465 -724 -1465 1 gnd
rlabel metal1 -639 -1367 -639 -1367 5 vdd
rlabel metal1 -634 -1455 -634 -1455 8 gnd
rlabel metal1 -676 -1367 -676 -1367 5 vdd
rlabel metal1 -671 -1455 -671 -1455 8 gnd
rlabel metal1 -767 -1758 -767 -1758 8 gnd
rlabel metal1 -730 -1758 -730 -1758 8 gnd
rlabel metal1 -820 -1768 -820 -1768 1 gnd
rlabel metal1 -735 -1670 -735 -1670 5 vdd
rlabel metal1 -772 -1670 -772 -1670 5 vdd
rlabel metal1 -768 -1640 -768 -1640 8 gnd
rlabel metal1 -773 -1552 -773 -1552 5 vdd
rlabel metal1 -731 -1640 -731 -1640 8 gnd
rlabel metal1 -736 -1552 -736 -1552 5 vdd
rlabel metal1 -821 -1650 -821 -1650 1 gnd
rlabel metal1 -660 -1660 -660 -1660 1 gnd
rlabel metal1 -575 -1562 -575 -1562 5 vdd
rlabel metal1 -570 -1650 -570 -1650 8 gnd
rlabel metal1 -612 -1562 -612 -1562 5 vdd
rlabel metal1 -607 -1650 -607 -1650 8 gnd
rlabel metal1 -929 -1894 -929 -1894 8 gnd
rlabel metal1 -934 -1806 -934 -1806 5 vdd
rlabel metal1 -892 -1894 -892 -1894 8 gnd
rlabel metal1 -897 -1806 -897 -1806 5 vdd
rlabel metal1 -982 -1904 -982 -1904 1 gnd
rlabel metal1 -867 -2007 -867 -2007 8 gnd
rlabel metal1 -872 -1919 -872 -1919 5 vdd
rlabel metal1 -1008 -1967 -1008 -1967 2 gnd
rlabel metal1 -920 -1962 -920 -1962 7 vdd
rlabel metal1 -920 -2002 -920 -2002 7 vdd
rlabel metal1 -1008 -2007 -1008 -2007 2 gnd
rlabel metal1 -640 -1944 -640 -1944 1 vdd
rlabel metal1 -552 -1888 -552 -1888 5 vdd
rlabel metal1 -547 -1976 -547 -1976 8 gnd
rlabel metal1 -589 -1888 -589 -1888 5 vdd
rlabel metal1 -584 -1976 -584 -1976 8 gnd
rlabel metal1 -736 -2008 -736 -2008 8 gnd
rlabel metal1 -741 -1920 -741 -1920 5 vdd
rlabel metal1 -699 -2008 -699 -2008 8 gnd
rlabel metal1 -704 -1920 -704 -1920 5 vdd
rlabel metal1 -789 -2018 -789 -2018 1 gnd
rlabel metal1 -546 -2166 -546 -2166 8 gnd
rlabel metal1 -551 -2078 -551 -2078 5 vdd
rlabel metal1 -509 -2166 -509 -2166 8 gnd
rlabel metal1 -514 -2078 -514 -2078 5 vdd
rlabel metal1 -602 -2134 -602 -2134 1 vdd
rlabel metal1 -822 -2816 -822 -2816 8 gnd
rlabel metal1 -827 -2728 -827 -2728 5 vdd
rlabel metal1 -785 -2816 -785 -2816 8 gnd
rlabel metal1 -790 -2728 -790 -2728 5 vdd
rlabel metal1 -875 -2826 -875 -2826 1 gnd
rlabel metal1 -1036 -2816 -1036 -2816 1 gnd
rlabel metal1 -951 -2718 -951 -2718 5 vdd
rlabel metal1 -946 -2806 -946 -2806 8 gnd
rlabel metal1 -988 -2718 -988 -2718 5 vdd
rlabel metal1 -983 -2806 -983 -2806 8 gnd
rlabel metal1 -675 -2710 -675 -2710 8 gnd
rlabel metal1 -680 -2622 -680 -2622 5 vdd
rlabel metal1 -638 -2710 -638 -2710 8 gnd
rlabel metal1 -643 -2622 -643 -2622 5 vdd
rlabel metal1 -728 -2720 -728 -2720 1 gnd
rlabel metal1 -853 -2689 -853 -2689 1 gnd
rlabel metal1 -768 -2591 -768 -2591 5 vdd
rlabel metal1 -763 -2679 -763 -2679 8 gnd
rlabel metal1 -805 -2591 -805 -2591 5 vdd
rlabel metal1 -800 -2679 -800 -2679 8 gnd
rlabel metal1 -688 -2193 -688 -2193 8 gnd
rlabel metal1 -693 -2105 -693 -2105 5 vdd
rlabel metal1 -651 -2193 -651 -2193 8 gnd
rlabel metal1 -656 -2105 -656 -2105 5 vdd
rlabel metal1 -744 -2161 -744 -2161 1 vdd
rlabel metal1 -1001 -2550 -1001 -2550 8 gnd
rlabel metal1 -964 -2550 -964 -2550 8 gnd
rlabel metal1 -1054 -2560 -1054 -2560 1 gnd
rlabel metal1 -969 -2462 -969 -2462 5 vdd
rlabel metal1 -1006 -2462 -1006 -2462 5 vdd
rlabel metal1 -1002 -2432 -1002 -2432 8 gnd
rlabel metal1 -1007 -2344 -1007 -2344 5 vdd
rlabel metal1 -965 -2432 -965 -2432 8 gnd
rlabel metal1 -970 -2344 -970 -2344 5 vdd
rlabel metal1 -1055 -2442 -1055 -2442 1 gnd
rlabel metal1 -894 -2452 -894 -2452 1 gnd
rlabel metal1 -809 -2354 -809 -2354 5 vdd
rlabel metal1 -804 -2442 -804 -2442 8 gnd
rlabel metal1 -846 -2354 -846 -2354 5 vdd
rlabel metal1 -841 -2442 -841 -2442 8 gnd
rlabel metal1 -1057 -2300 -1057 -2300 8 gnd
rlabel metal1 -1062 -2212 -1062 -2212 5 vdd
rlabel metal1 -1020 -2300 -1020 -2300 8 gnd
rlabel metal1 -1025 -2212 -1025 -2212 5 vdd
rlabel metal1 -1110 -2310 -1110 -2310 1 gnd
rlabel metal1 -949 -2320 -949 -2320 1 gnd
rlabel metal1 -864 -2222 -864 -2222 5 vdd
rlabel metal1 -859 -2310 -859 -2310 8 gnd
rlabel metal1 -901 -2222 -901 -2222 5 vdd
rlabel metal1 -896 -2310 -896 -2310 8 gnd
rlabel metal1 -958 -377 -958 -377 1 a0
rlabel metal1 -966 -407 -966 -406 1 b0
rlabel metal1 -965 -648 -965 -648 1 a1
rlabel metal1 -976 -678 -976 -678 1 b1
rlabel metal1 -968 -1080 -968 -1080 1 a2
rlabel metal1 -976 -1110 -976 -1110 1 b2
rlabel metal1 -1030 -1831 -1030 -1831 1 a3
rlabel metal1 -1039 -1862 -1039 -1862 1 b3
rlabel metal1 -1289 -249 -1289 -249 1 c0
rlabel metal1 -1289 -291 -1289 -291 1 p0
rlabel metal1 -390 -504 -390 -504 1 c1
rlabel metal1 -389 -546 -389 -546 1 p1
rlabel metal1 -223 -776 -223 -776 1 c2
rlabel metal1 -210 -817 -210 -817 1 p2
rlabel metal1 -209 -1207 -209 -1207 1 c3
rlabel metal1 -203 -1248 -203 -1248 1 p3
rlabel metal1 -71 -1241 -71 -1241 1 s3
rlabel metal1 -68 -811 -68 -811 1 s2
rlabel metal1 -254 -539 -254 -539 1 s1
rlabel metal1 -265 -286 -265 -286 1 s0
rlabel metal1 -810 -408 -810 -408 1 g0
rlabel metal1 -817 -680 -817 -680 1 g1
rlabel metal1 -813 -1111 -813 -1111 1 g2
rlabel metal1 -872 -1862 -872 -1862 1 g3
rlabel metal1 -409 -2007 -409 -2007 8 gnd
rlabel metal1 -414 -1919 -414 -1919 5 vdd
rlabel metal1 -372 -2007 -372 -2007 8 gnd
rlabel metal1 -377 -1919 -377 -1919 5 vdd
rlabel metal1 -465 -1975 -465 -1975 1 vdd
rlabel metal1 -361 -1975 -361 -1975 1 cout
<< end >>
